package Step;
import Operation::*;
import Types::*;
import Vector::*;
import FShow::*;
import Debug::*;
import PMU::*;
import RamulatorArbiter::*;
import RandomLoad::*;

(* synthesize *)
module mkHypernode_6034 (Operation_IFC);
    Operation_IFC mod_1_inner <- mkReshape(2, 64);
    Operation_IFC mod_1 <- mkDebugOperation(mod_1_inner, "mod_1");
    Operation_IFC mod_2_inner <- mkFlatten(1);
    Operation_IFC mod_2 <- mkDebugOperation(mod_2_inner, "mod_2");
    Operation_IFC mod_3_inner <- mkFlatten(2);
    Operation_IFC mod_3 <- mkDebugOperation(mod_3_inner, "mod_3");
    Operation_IFC mod_4_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4 <- mkDebugOperation(mod_4_inner, "mod_4");
    Broadcast_IFC#(4) mod_5_inner <- mkBroadcast(4);
    Operation_IFC mod_5 <- mkDebugOperation(mod_5_inner.op, "mod_5");
    PMU_IFC mod_6_bufferize <- mkPMU(2);
    Operation_IFC mod_6_inner = mod_6_bufferize.operation;
    Operation_IFC mod_6 <- mkDebugOperation(mod_6_inner, "mod_6");
    Broadcast_IFC#(2) mod_7_inner <- mkBroadcast(2);
    Operation_IFC mod_7 <- mkDebugOperation(mod_7_inner.op, "mod_7");
    PMU_IFC mod_8_bufferize <- mkPMU(1);
    Operation_IFC mod_8_inner = mod_8_bufferize.operation;
    Operation_IFC mod_8 <- mkDebugOperation(mod_8_inner, "mod_8");
    Operation_IFC mod_9_inner <- mkBinaryMap(1156, matmul_t_tile);
    Operation_IFC mod_9 <- mkDebugOperation(mod_9_inner, "mod_9");
    Operation_IFC mod_10_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_10 <- mkDebugOperation(mod_10_inner, "mod_10");
    Operation_IFC mod_11_inner <- mkBinaryMap(1924, mul_tile);
    Operation_IFC mod_11 <- mkDebugOperation(mod_11_inner, "mod_11");
    PMU_IFC mod_12_bufferize <- mkPMU(1);
    Operation_IFC mod_12_inner = mod_12_bufferize.operation;
    Operation_IFC mod_12 <- mkDebugOperation(mod_12_inner, "mod_12");
    Operation_IFC mod_13_inner <- mkBinaryMap(2563, matmul_t_tile);
    Operation_IFC mod_13 <- mkDebugOperation(mod_13_inner, "mod_13");
    Operation_IFC mod_14_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_14 <- mkDebugOperation(mod_14_inner, "mod_14");
    Operation_IFC mod_15_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_15 <- mkDebugOperation(mod_15_inner, "mod_15");
    Operation_IFC mod_16_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_16 <- mkDebugOperation(mod_16_inner, "mod_16");
    Operation_IFC mod_17_inner <- mkBinaryMap(2823, mul_tile);
    Operation_IFC mod_17 <- mkDebugOperation(mod_17_inner, "mod_17");
    PMU_IFC mod_18_bufferize <- mkPMU(1);
    Operation_IFC mod_18_inner = mod_18_bufferize.operation;
    Operation_IFC mod_18 <- mkDebugOperation(mod_18_inner, "mod_18");
    PMU_IFC mod_19_bufferize <- mkPMU(2);
    Operation_IFC mod_19_inner = mod_19_bufferize.operation;
    Operation_IFC mod_19 <- mkDebugOperation(mod_19_inner, "mod_19");
    PMU_IFC mod_20_bufferize <- mkPMU(2);
    Operation_IFC mod_20_inner = mod_20_bufferize.operation;
    Operation_IFC mod_20 <- mkDebugOperation(mod_20_inner, "mod_20");
    Operation_IFC mod_21_inner <- mkRepeatStatic(8);
    Operation_IFC mod_21 <- mkDebugOperation(mod_21_inner, "mod_21");
    Operation_IFC mod_22_inner <- mkFlatten(1);
    Operation_IFC mod_22 <- mkDebugOperation(mod_22_inner, "mod_22");
    Operation_IFC mod_23_inner <- mkFlatten(0);
    Operation_IFC mod_23 <- mkDebugOperation(mod_23_inner, "mod_23");
    Operation_IFC mod_24_inner <- mkRepeatStatic(3);
    Operation_IFC mod_24 <- mkDebugOperation(mod_24_inner, "mod_24");
    Operation_IFC mod_25_inner <- mkUnaryMap(1796, silu_tile);
    Operation_IFC mod_25 <- mkDebugOperation(mod_25_inner, "mod_25");
    Operation_IFC mod_26_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_26 <- mkDebugOperation(mod_26_inner, "mod_26");
    Operation_IFC mod_27_inner <- mkBinaryMap(1668, matmul_t_tile);
    Operation_IFC mod_27 <- mkDebugOperation(mod_27_inner, "mod_27");
    PMU_IFC mod_28_bufferize <- mkPMU(2);
    Operation_IFC mod_28_inner = mod_28_bufferize.operation;
    Operation_IFC mod_28 <- mkDebugOperation(mod_28_inner, "mod_28");
    Operation_IFC mod_29_inner <- mkRepeatStatic(8);
    Operation_IFC mod_29 <- mkDebugOperation(mod_29_inner, "mod_29");
    Operation_IFC mod_30_inner <- mkFlatten(1);
    Operation_IFC mod_30 <- mkDebugOperation(mod_30_inner, "mod_30");
    Operation_IFC mod_31_inner <- mkFlatten(0);
    Operation_IFC mod_31 <- mkDebugOperation(mod_31_inner, "mod_31");
    PMU_IFC mod_32_bufferize <- mkPMU(1);
    Operation_IFC mod_32_inner = mod_32_bufferize.operation;
    Operation_IFC mod_32 <- mkDebugOperation(mod_32_inner, "mod_32");
    Operation_IFC mod_33_inner <- mkRepeatStatic(16);
    Operation_IFC mod_33 <- mkDebugOperation(mod_33_inner, "mod_33");
    PMU_IFC mod_34_bufferize <- mkPMU(2);
    Operation_IFC mod_34_inner = mod_34_bufferize.operation;
    Operation_IFC mod_34 <- mkDebugOperation(mod_34_inner, "mod_34");
    Operation_IFC mod_35_inner <- mkRepeatStatic(8);
    Operation_IFC mod_35 <- mkDebugOperation(mod_35_inner, "mod_35");
    Operation_IFC mod_36_inner <- mkFlatten(1);
    Operation_IFC mod_36 <- mkDebugOperation(mod_36_inner, "mod_36");
    Operation_IFC mod_37_inner <- mkFlatten(0);
    Operation_IFC mod_37 <- mkDebugOperation(mod_37_inner, "mod_37");
    Operation_IFC mod_38_inner <- mkRepeatStatic(16);
    Operation_IFC mod_38 <- mkDebugOperation(mod_38_inner, "mod_38");
    Operation_IFC mod_39_inner <- mkRepeatStatic(2);
    Operation_IFC mod_39 <- mkDebugOperation(mod_39_inner, "mod_39");
    PMU_IFC mod_40_bufferize <- mkPMU(2);
    Operation_IFC mod_40_inner = mod_40_bufferize.operation;
    Operation_IFC mod_40 <- mkDebugOperation(mod_40_inner, "mod_40");
    rule rule_1;
        ChannelMessage t;
        t <- mod_28.get(1);
        mod_27.put(1, t);
    endrule
    rule rule_2;
        ChannelMessage t;
        t <- mod_10.get(0);
        mod_11.put(0, t);
    endrule
    rule rule_3;
        ChannelMessage t;
        t <- mod_15.get(0);
        mod_19.put(0, t);
    endrule
    rule rule_4;
        ChannelMessage t;
        t <- mod_28.get(0);
        mod_29.put(0, t);
    endrule
    rule rule_5;
        ChannelMessage t;
        t <- mod_4.get(1);
        mod_5.put(0, t);
    endrule
    rule rule_6;
        ChannelMessage t;
        t <- mod_16.get(0);
        mod_18.put(0, t);
    endrule
    rule rule_7;
        ChannelMessage t;
        t <- mod_14.get(0);
        mod_15.put(0, t);
    endrule
    rule rule_8;
        ChannelMessage t;
        t <- mod_30.get(0);
        mod_28.put(0, t);
    endrule
    rule rule_9;
        ChannelMessage t;
        t <- mod_33.get(0);
        mod_32.put(1, t);
    endrule
    rule rule_10;
        ChannelMessage t;
        t <- mod_8.get(1);
        mod_9.put(0, t);
    endrule
    rule rule_11;
        ChannelMessage t;
        t <- mod_34.get(0);
        mod_35.put(0, t);
    endrule
    rule rule_12;
        ChannelMessage t;
        t <- mod_40.get(1);
        mod_4.put(1, t);
    endrule
    rule rule_13;
        ChannelMessage t;
        t <- mod_25.get(0);
        mod_11.put(1, t);
    endrule
    rule rule_14;
        ChannelMessage t;
        t <- mod_23.get(0);
        mod_22.put(0, t);
    endrule
    rule rule_15;
        ChannelMessage t;
        t <- mod_20.get(0);
        mod_21.put(0, t);
    endrule
    rule rule_16;
        ChannelMessage t;
        t <- mod_18.get(0);
        mod_18.put(1, t);
    endrule
    rule rule_17;
        ChannelMessage t;
        t <- mod_20.get(1);
        mod_13.put(1, t);
    endrule
    rule rule_18;
        ChannelMessage t;
        t <- mod_18.get(1);
        mod_16.put(1, t);
    endrule
    rule rule_19;
        ChannelMessage t;
        t <- mod_29.get(0);
        mod_28.put(1, t);
    endrule
    rule rule_20;
        ChannelMessage t;
        t <- mod_34.get(1);
        mod_9.put(1, t);
    endrule
    rule rule_21;
        ChannelMessage t;
        t <- mod_32.get(1);
        mod_27.put(0, t);
    endrule
    rule rule_22;
        ChannelMessage t;
        t <- mod_40.get(0);
        mod_40.put(1, t);
    endrule
    rule rule_23;
        ChannelMessage t;
        t <- mod_32.get(0);
        mod_33.put(0, t);
    endrule
    rule rule_24;
        ChannelMessage t;
        t <- mod_12.get(1);
        mod_13.put(0, t);
    endrule
    rule rule_25;
        ChannelMessage t;
        t <- mod_24.get(0);
        mod_12.put(1, t);
    endrule
    rule rule_26;
        ChannelMessage t;
        t <- mod_21.get(0);
        mod_20.put(1, t);
    endrule
    rule rule_27;
        ChannelMessage t;
        t <- mod_13.get(0);
        mod_14.put(0, t);
    endrule
    rule rule_28;
        ChannelMessage t;
        t <- mod_2.get(0);
        mod_3.put(0, t);
    endrule
    rule rule_29;
        ChannelMessage t;
        t <- mod_19.get(1);
        mod_15.put(1, t);
    endrule
    rule rule_30;
        ChannelMessage t;
        t <- mod_26.get(0);
        mod_25.put(0, t);
    endrule
    rule rule_31;
        ChannelMessage t;
        t <- mod_35.get(0);
        mod_34.put(1, t);
    endrule
    rule rule_32;
        ChannelMessage t;
        t <- mod_7.get(0);
        mod_32.put(0, t);
    endrule
    rule rule_33;
        ChannelMessage t;
        t <- mod_6.get(0);
        mod_39.put(0, t);
    endrule
    rule rule_34;
        ChannelMessage t;
        t <- mod_7.get(1);
        mod_8.put(0, t);
    endrule
    rule rule_35;
        ChannelMessage t;
        t <- mod_8.get(0);
        mod_38.put(0, t);
    endrule
    rule rule_36;
        ChannelMessage t;
        t <- mod_31.get(0);
        mod_30.put(0, t);
    endrule
    rule rule_37;
        ChannelMessage t;
        t <- mod_16.get(1);
        mod_17.put(1, t);
    endrule
    rule rule_38;
        ChannelMessage t;
        t <- mod_11.get(0);
        mod_12.put(0, t);
    endrule
    rule rule_39;
        ChannelMessage t;
        t <- mod_1.get(0);
        mod_2.put(0, t);
    endrule
    rule rule_40;
        ChannelMessage t;
        t <- mod_38.get(0);
        mod_8.put(1, t);
    endrule
    rule rule_41;
        ChannelMessage t;
        t <- mod_6.get(1);
        mod_7.put(0, t);
    endrule
    rule rule_42;
        ChannelMessage t;
        t <- mod_5.get(3);
        mod_6.put(0, t);
    endrule
    rule rule_43;
        ChannelMessage t;
        t <- mod_36.get(0);
        mod_34.put(0, t);
    endrule
    rule rule_44;
        ChannelMessage t;
        t <- mod_19.get(0);
        mod_19.put(1, t);
    endrule
    rule rule_45;
        ChannelMessage t;
        t <- mod_22.get(0);
        mod_20.put(0, t);
    endrule
    rule rule_46;
        ChannelMessage t;
        t <- mod_15.get(1);
        mod_16.put(0, t);
    endrule
    rule rule_47;
        ChannelMessage t;
        t <- mod_37.get(0);
        mod_36.put(0, t);
    endrule
    rule rule_48;
        ChannelMessage t;
        t <- mod_27.get(0);
        mod_26.put(0, t);
    endrule
    rule rule_49;
        ChannelMessage t;
        t <- mod_39.get(0);
        mod_6.put(1, t);
    endrule
    rule rule_50;
        ChannelMessage t;
        t <- mod_3.get(0);
        mod_4.put(0, t);
    endrule
    rule rule_51;
        ChannelMessage t;
        t <- mod_9.get(0);
        mod_10.put(0, t);
    endrule
    rule rule_52;
        ChannelMessage t;
        t <- mod_4.get(0);
        mod_40.put(0, t);
    endrule
    rule rule_53;
        ChannelMessage t;
        t <- mod_12.get(0);
        mod_24.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1.put(0, t);
        end
        if (i == 1) begin
            mod_17.put(0, t);
        end
        if (i == 2) begin
            mod_23.put(0, t);
        end
        if (i == 3) begin
            mod_31.put(0, t);
        end
        if (i == 4) begin
            mod_37.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_5.get(0);
        end
        if (i == 2) begin
            t <- mod_5.get(1);
        end
        if (i == 1) begin
            t <- mod_5.get(2);
        end
        if (i == 0) begin
            t <- mod_17.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6035 (Operation_IFC);
    Operation_IFC mod_42_inner <- mkReshape(2, 64);
    Operation_IFC mod_42 <- mkDebugOperation(mod_42_inner, "mod_42");
    Operation_IFC mod_43_inner <- mkFlatten(1);
    Operation_IFC mod_43 <- mkDebugOperation(mod_43_inner, "mod_43");
    Operation_IFC mod_44_inner <- mkFlatten(2);
    Operation_IFC mod_44 <- mkDebugOperation(mod_44_inner, "mod_44");
    Operation_IFC mod_45_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_45 <- mkDebugOperation(mod_45_inner, "mod_45");
    Broadcast_IFC#(4) mod_46_inner <- mkBroadcast(4);
    Operation_IFC mod_46 <- mkDebugOperation(mod_46_inner.op, "mod_46");
    PMU_IFC mod_47_bufferize <- mkPMU(2);
    Operation_IFC mod_47_inner = mod_47_bufferize.operation;
    Operation_IFC mod_47 <- mkDebugOperation(mod_47_inner, "mod_47");
    Broadcast_IFC#(2) mod_48_inner <- mkBroadcast(2);
    Operation_IFC mod_48 <- mkDebugOperation(mod_48_inner.op, "mod_48");
    PMU_IFC mod_49_bufferize <- mkPMU(1);
    Operation_IFC mod_49_inner = mod_49_bufferize.operation;
    Operation_IFC mod_49 <- mkDebugOperation(mod_49_inner, "mod_49");
    Operation_IFC mod_50_inner <- mkBinaryMap(1155, matmul_t_tile);
    Operation_IFC mod_50 <- mkDebugOperation(mod_50_inner, "mod_50");
    Operation_IFC mod_51_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_51 <- mkDebugOperation(mod_51_inner, "mod_51");
    Operation_IFC mod_52_inner <- mkBinaryMap(1923, mul_tile);
    Operation_IFC mod_52 <- mkDebugOperation(mod_52_inner, "mod_52");
    PMU_IFC mod_53_bufferize <- mkPMU(1);
    Operation_IFC mod_53_inner = mod_53_bufferize.operation;
    Operation_IFC mod_53 <- mkDebugOperation(mod_53_inner, "mod_53");
    Operation_IFC mod_54_inner <- mkBinaryMap(2561, matmul_t_tile);
    Operation_IFC mod_54 <- mkDebugOperation(mod_54_inner, "mod_54");
    Operation_IFC mod_55_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_55 <- mkDebugOperation(mod_55_inner, "mod_55");
    Operation_IFC mod_56_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_56 <- mkDebugOperation(mod_56_inner, "mod_56");
    Operation_IFC mod_57_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_57 <- mkDebugOperation(mod_57_inner, "mod_57");
    Operation_IFC mod_58_inner <- mkBinaryMap(2822, mul_tile);
    Operation_IFC mod_58 <- mkDebugOperation(mod_58_inner, "mod_58");
    PMU_IFC mod_59_bufferize <- mkPMU(1);
    Operation_IFC mod_59_inner = mod_59_bufferize.operation;
    Operation_IFC mod_59 <- mkDebugOperation(mod_59_inner, "mod_59");
    PMU_IFC mod_60_bufferize <- mkPMU(2);
    Operation_IFC mod_60_inner = mod_60_bufferize.operation;
    Operation_IFC mod_60 <- mkDebugOperation(mod_60_inner, "mod_60");
    PMU_IFC mod_61_bufferize <- mkPMU(2);
    Operation_IFC mod_61_inner = mod_61_bufferize.operation;
    Operation_IFC mod_61 <- mkDebugOperation(mod_61_inner, "mod_61");
    Operation_IFC mod_62_inner <- mkRepeatStatic(8);
    Operation_IFC mod_62 <- mkDebugOperation(mod_62_inner, "mod_62");
    Operation_IFC mod_63_inner <- mkFlatten(1);
    Operation_IFC mod_63 <- mkDebugOperation(mod_63_inner, "mod_63");
    Operation_IFC mod_64_inner <- mkFlatten(0);
    Operation_IFC mod_64 <- mkDebugOperation(mod_64_inner, "mod_64");
    Operation_IFC mod_65_inner <- mkRepeatStatic(3);
    Operation_IFC mod_65 <- mkDebugOperation(mod_65_inner, "mod_65");
    Operation_IFC mod_66_inner <- mkUnaryMap(1795, silu_tile);
    Operation_IFC mod_66 <- mkDebugOperation(mod_66_inner, "mod_66");
    Operation_IFC mod_67_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_67 <- mkDebugOperation(mod_67_inner, "mod_67");
    Operation_IFC mod_68_inner <- mkBinaryMap(1667, matmul_t_tile);
    Operation_IFC mod_68 <- mkDebugOperation(mod_68_inner, "mod_68");
    PMU_IFC mod_69_bufferize <- mkPMU(2);
    Operation_IFC mod_69_inner = mod_69_bufferize.operation;
    Operation_IFC mod_69 <- mkDebugOperation(mod_69_inner, "mod_69");
    Operation_IFC mod_70_inner <- mkRepeatStatic(8);
    Operation_IFC mod_70 <- mkDebugOperation(mod_70_inner, "mod_70");
    Operation_IFC mod_71_inner <- mkFlatten(1);
    Operation_IFC mod_71 <- mkDebugOperation(mod_71_inner, "mod_71");
    Operation_IFC mod_72_inner <- mkFlatten(0);
    Operation_IFC mod_72 <- mkDebugOperation(mod_72_inner, "mod_72");
    PMU_IFC mod_73_bufferize <- mkPMU(1);
    Operation_IFC mod_73_inner = mod_73_bufferize.operation;
    Operation_IFC mod_73 <- mkDebugOperation(mod_73_inner, "mod_73");
    Operation_IFC mod_74_inner <- mkRepeatStatic(16);
    Operation_IFC mod_74 <- mkDebugOperation(mod_74_inner, "mod_74");
    PMU_IFC mod_75_bufferize <- mkPMU(2);
    Operation_IFC mod_75_inner = mod_75_bufferize.operation;
    Operation_IFC mod_75 <- mkDebugOperation(mod_75_inner, "mod_75");
    Operation_IFC mod_76_inner <- mkRepeatStatic(8);
    Operation_IFC mod_76 <- mkDebugOperation(mod_76_inner, "mod_76");
    Operation_IFC mod_77_inner <- mkFlatten(1);
    Operation_IFC mod_77 <- mkDebugOperation(mod_77_inner, "mod_77");
    Operation_IFC mod_78_inner <- mkFlatten(0);
    Operation_IFC mod_78 <- mkDebugOperation(mod_78_inner, "mod_78");
    Operation_IFC mod_79_inner <- mkRepeatStatic(16);
    Operation_IFC mod_79 <- mkDebugOperation(mod_79_inner, "mod_79");
    Operation_IFC mod_80_inner <- mkRepeatStatic(2);
    Operation_IFC mod_80 <- mkDebugOperation(mod_80_inner, "mod_80");
    PMU_IFC mod_81_bufferize <- mkPMU(2);
    Operation_IFC mod_81_inner = mod_81_bufferize.operation;
    Operation_IFC mod_81 <- mkDebugOperation(mod_81_inner, "mod_81");
    rule rule_54;
        ChannelMessage t;
        t <- mod_60.get(0);
        mod_60.put(1, t);
    endrule
    rule rule_55;
        ChannelMessage t;
        t <- mod_73.get(1);
        mod_68.put(0, t);
    endrule
    rule rule_56;
        ChannelMessage t;
        t <- mod_48.get(0);
        mod_73.put(0, t);
    endrule
    rule rule_57;
        ChannelMessage t;
        t <- mod_53.get(1);
        mod_54.put(0, t);
    endrule
    rule rule_58;
        ChannelMessage t;
        t <- mod_79.get(0);
        mod_49.put(1, t);
    endrule
    rule rule_59;
        ChannelMessage t;
        t <- mod_47.get(1);
        mod_48.put(0, t);
    endrule
    rule rule_60;
        ChannelMessage t;
        t <- mod_76.get(0);
        mod_75.put(1, t);
    endrule
    rule rule_61;
        ChannelMessage t;
        t <- mod_69.get(0);
        mod_70.put(0, t);
    endrule
    rule rule_62;
        ChannelMessage t;
        t <- mod_70.get(0);
        mod_69.put(1, t);
    endrule
    rule rule_63;
        ChannelMessage t;
        t <- mod_65.get(0);
        mod_53.put(1, t);
    endrule
    rule rule_64;
        ChannelMessage t;
        t <- mod_61.get(0);
        mod_62.put(0, t);
    endrule
    rule rule_65;
        ChannelMessage t;
        t <- mod_47.get(0);
        mod_80.put(0, t);
    endrule
    rule rule_66;
        ChannelMessage t;
        t <- mod_72.get(0);
        mod_71.put(0, t);
    endrule
    rule rule_67;
        ChannelMessage t;
        t <- mod_74.get(0);
        mod_73.put(1, t);
    endrule
    rule rule_68;
        ChannelMessage t;
        t <- mod_81.get(1);
        mod_45.put(1, t);
    endrule
    rule rule_69;
        ChannelMessage t;
        t <- mod_49.get(1);
        mod_50.put(0, t);
    endrule
    rule rule_70;
        ChannelMessage t;
        t <- mod_52.get(0);
        mod_53.put(0, t);
    endrule
    rule rule_71;
        ChannelMessage t;
        t <- mod_60.get(1);
        mod_56.put(1, t);
    endrule
    rule rule_72;
        ChannelMessage t;
        t <- mod_75.get(0);
        mod_76.put(0, t);
    endrule
    rule rule_73;
        ChannelMessage t;
        t <- mod_57.get(0);
        mod_59.put(0, t);
    endrule
    rule rule_74;
        ChannelMessage t;
        t <- mod_57.get(1);
        mod_58.put(1, t);
    endrule
    rule rule_75;
        ChannelMessage t;
        t <- mod_42.get(0);
        mod_43.put(0, t);
    endrule
    rule rule_76;
        ChannelMessage t;
        t <- mod_53.get(0);
        mod_65.put(0, t);
    endrule
    rule rule_77;
        ChannelMessage t;
        t <- mod_54.get(0);
        mod_55.put(0, t);
    endrule
    rule rule_78;
        ChannelMessage t;
        t <- mod_56.get(1);
        mod_57.put(0, t);
    endrule
    rule rule_79;
        ChannelMessage t;
        t <- mod_59.get(0);
        mod_59.put(1, t);
    endrule
    rule rule_80;
        ChannelMessage t;
        t <- mod_69.get(1);
        mod_68.put(1, t);
    endrule
    rule rule_81;
        ChannelMessage t;
        t <- mod_46.get(3);
        mod_47.put(0, t);
    endrule
    rule rule_82;
        ChannelMessage t;
        t <- mod_71.get(0);
        mod_69.put(0, t);
    endrule
    rule rule_83;
        ChannelMessage t;
        t <- mod_75.get(1);
        mod_50.put(1, t);
    endrule
    rule rule_84;
        ChannelMessage t;
        t <- mod_77.get(0);
        mod_75.put(0, t);
    endrule
    rule rule_85;
        ChannelMessage t;
        t <- mod_45.get(0);
        mod_81.put(0, t);
    endrule
    rule rule_86;
        ChannelMessage t;
        t <- mod_61.get(1);
        mod_54.put(1, t);
    endrule
    rule rule_87;
        ChannelMessage t;
        t <- mod_48.get(1);
        mod_49.put(0, t);
    endrule
    rule rule_88;
        ChannelMessage t;
        t <- mod_45.get(1);
        mod_46.put(0, t);
    endrule
    rule rule_89;
        ChannelMessage t;
        t <- mod_43.get(0);
        mod_44.put(0, t);
    endrule
    rule rule_90;
        ChannelMessage t;
        t <- mod_67.get(0);
        mod_66.put(0, t);
    endrule
    rule rule_91;
        ChannelMessage t;
        t <- mod_78.get(0);
        mod_77.put(0, t);
    endrule
    rule rule_92;
        ChannelMessage t;
        t <- mod_55.get(0);
        mod_56.put(0, t);
    endrule
    rule rule_93;
        ChannelMessage t;
        t <- mod_64.get(0);
        mod_63.put(0, t);
    endrule
    rule rule_94;
        ChannelMessage t;
        t <- mod_68.get(0);
        mod_67.put(0, t);
    endrule
    rule rule_95;
        ChannelMessage t;
        t <- mod_49.get(0);
        mod_79.put(0, t);
    endrule
    rule rule_96;
        ChannelMessage t;
        t <- mod_81.get(0);
        mod_81.put(1, t);
    endrule
    rule rule_97;
        ChannelMessage t;
        t <- mod_63.get(0);
        mod_61.put(0, t);
    endrule
    rule rule_98;
        ChannelMessage t;
        t <- mod_59.get(1);
        mod_57.put(1, t);
    endrule
    rule rule_99;
        ChannelMessage t;
        t <- mod_56.get(0);
        mod_60.put(0, t);
    endrule
    rule rule_100;
        ChannelMessage t;
        t <- mod_66.get(0);
        mod_52.put(1, t);
    endrule
    rule rule_101;
        ChannelMessage t;
        t <- mod_51.get(0);
        mod_52.put(0, t);
    endrule
    rule rule_102;
        ChannelMessage t;
        t <- mod_80.get(0);
        mod_47.put(1, t);
    endrule
    rule rule_103;
        ChannelMessage t;
        t <- mod_44.get(0);
        mod_45.put(0, t);
    endrule
    rule rule_104;
        ChannelMessage t;
        t <- mod_50.get(0);
        mod_51.put(0, t);
    endrule
    rule rule_105;
        ChannelMessage t;
        t <- mod_62.get(0);
        mod_61.put(1, t);
    endrule
    rule rule_106;
        ChannelMessage t;
        t <- mod_73.get(0);
        mod_74.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_42.put(0, t);
        end
        if (i == 1) begin
            mod_58.put(0, t);
        end
        if (i == 2) begin
            mod_64.put(0, t);
        end
        if (i == 3) begin
            mod_72.put(0, t);
        end
        if (i == 4) begin
            mod_78.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 2) begin
            t <- mod_46.get(0);
        end
        if (i == 1) begin
            t <- mod_46.get(1);
        end
        if (i == 3) begin
            t <- mod_46.get(2);
        end
        if (i == 0) begin
            t <- mod_58.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6036 (Operation_IFC);
    Operation_IFC mod_83_inner <- mkReshape(2, 64);
    Operation_IFC mod_83 <- mkDebugOperation(mod_83_inner, "mod_83");
    Operation_IFC mod_84_inner <- mkFlatten(1);
    Operation_IFC mod_84 <- mkDebugOperation(mod_84_inner, "mod_84");
    Operation_IFC mod_85_inner <- mkFlatten(2);
    Operation_IFC mod_85 <- mkDebugOperation(mod_85_inner, "mod_85");
    Operation_IFC mod_86_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_86 <- mkDebugOperation(mod_86_inner, "mod_86");
    Broadcast_IFC#(4) mod_87_inner <- mkBroadcast(4);
    Operation_IFC mod_87 <- mkDebugOperation(mod_87_inner.op, "mod_87");
    PMU_IFC mod_88_bufferize <- mkPMU(2);
    Operation_IFC mod_88_inner = mod_88_bufferize.operation;
    Operation_IFC mod_88 <- mkDebugOperation(mod_88_inner, "mod_88");
    Broadcast_IFC#(2) mod_89_inner <- mkBroadcast(2);
    Operation_IFC mod_89 <- mkDebugOperation(mod_89_inner.op, "mod_89");
    PMU_IFC mod_90_bufferize <- mkPMU(1);
    Operation_IFC mod_90_inner = mod_90_bufferize.operation;
    Operation_IFC mod_90 <- mkDebugOperation(mod_90_inner, "mod_90");
    Operation_IFC mod_91_inner <- mkBinaryMap(1154, matmul_t_tile);
    Operation_IFC mod_91 <- mkDebugOperation(mod_91_inner, "mod_91");
    Operation_IFC mod_92_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_92 <- mkDebugOperation(mod_92_inner, "mod_92");
    Operation_IFC mod_93_inner <- mkBinaryMap(1922, mul_tile);
    Operation_IFC mod_93 <- mkDebugOperation(mod_93_inner, "mod_93");
    PMU_IFC mod_94_bufferize <- mkPMU(1);
    Operation_IFC mod_94_inner = mod_94_bufferize.operation;
    Operation_IFC mod_94 <- mkDebugOperation(mod_94_inner, "mod_94");
    Operation_IFC mod_95_inner <- mkBinaryMap(2559, matmul_t_tile);
    Operation_IFC mod_95 <- mkDebugOperation(mod_95_inner, "mod_95");
    Operation_IFC mod_96_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_96 <- mkDebugOperation(mod_96_inner, "mod_96");
    Operation_IFC mod_97_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_97 <- mkDebugOperation(mod_97_inner, "mod_97");
    Operation_IFC mod_98_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_98 <- mkDebugOperation(mod_98_inner, "mod_98");
    Operation_IFC mod_99_inner <- mkBinaryMap(2821, mul_tile);
    Operation_IFC mod_99 <- mkDebugOperation(mod_99_inner, "mod_99");
    PMU_IFC mod_100_bufferize <- mkPMU(1);
    Operation_IFC mod_100_inner = mod_100_bufferize.operation;
    Operation_IFC mod_100 <- mkDebugOperation(mod_100_inner, "mod_100");
    PMU_IFC mod_101_bufferize <- mkPMU(2);
    Operation_IFC mod_101_inner = mod_101_bufferize.operation;
    Operation_IFC mod_101 <- mkDebugOperation(mod_101_inner, "mod_101");
    PMU_IFC mod_102_bufferize <- mkPMU(2);
    Operation_IFC mod_102_inner = mod_102_bufferize.operation;
    Operation_IFC mod_102 <- mkDebugOperation(mod_102_inner, "mod_102");
    Operation_IFC mod_103_inner <- mkRepeatStatic(8);
    Operation_IFC mod_103 <- mkDebugOperation(mod_103_inner, "mod_103");
    Operation_IFC mod_104_inner <- mkFlatten(1);
    Operation_IFC mod_104 <- mkDebugOperation(mod_104_inner, "mod_104");
    Operation_IFC mod_105_inner <- mkFlatten(0);
    Operation_IFC mod_105 <- mkDebugOperation(mod_105_inner, "mod_105");
    Operation_IFC mod_106_inner <- mkRepeatStatic(3);
    Operation_IFC mod_106 <- mkDebugOperation(mod_106_inner, "mod_106");
    Operation_IFC mod_107_inner <- mkUnaryMap(1794, silu_tile);
    Operation_IFC mod_107 <- mkDebugOperation(mod_107_inner, "mod_107");
    Operation_IFC mod_108_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_108 <- mkDebugOperation(mod_108_inner, "mod_108");
    Operation_IFC mod_109_inner <- mkBinaryMap(1666, matmul_t_tile);
    Operation_IFC mod_109 <- mkDebugOperation(mod_109_inner, "mod_109");
    PMU_IFC mod_110_bufferize <- mkPMU(2);
    Operation_IFC mod_110_inner = mod_110_bufferize.operation;
    Operation_IFC mod_110 <- mkDebugOperation(mod_110_inner, "mod_110");
    Operation_IFC mod_111_inner <- mkRepeatStatic(8);
    Operation_IFC mod_111 <- mkDebugOperation(mod_111_inner, "mod_111");
    Operation_IFC mod_112_inner <- mkFlatten(1);
    Operation_IFC mod_112 <- mkDebugOperation(mod_112_inner, "mod_112");
    Operation_IFC mod_113_inner <- mkFlatten(0);
    Operation_IFC mod_113 <- mkDebugOperation(mod_113_inner, "mod_113");
    PMU_IFC mod_114_bufferize <- mkPMU(1);
    Operation_IFC mod_114_inner = mod_114_bufferize.operation;
    Operation_IFC mod_114 <- mkDebugOperation(mod_114_inner, "mod_114");
    Operation_IFC mod_115_inner <- mkRepeatStatic(16);
    Operation_IFC mod_115 <- mkDebugOperation(mod_115_inner, "mod_115");
    PMU_IFC mod_116_bufferize <- mkPMU(2);
    Operation_IFC mod_116_inner = mod_116_bufferize.operation;
    Operation_IFC mod_116 <- mkDebugOperation(mod_116_inner, "mod_116");
    Operation_IFC mod_117_inner <- mkRepeatStatic(8);
    Operation_IFC mod_117 <- mkDebugOperation(mod_117_inner, "mod_117");
    Operation_IFC mod_118_inner <- mkFlatten(1);
    Operation_IFC mod_118 <- mkDebugOperation(mod_118_inner, "mod_118");
    Operation_IFC mod_119_inner <- mkFlatten(0);
    Operation_IFC mod_119 <- mkDebugOperation(mod_119_inner, "mod_119");
    Operation_IFC mod_120_inner <- mkRepeatStatic(16);
    Operation_IFC mod_120 <- mkDebugOperation(mod_120_inner, "mod_120");
    Operation_IFC mod_121_inner <- mkRepeatStatic(2);
    Operation_IFC mod_121 <- mkDebugOperation(mod_121_inner, "mod_121");
    PMU_IFC mod_122_bufferize <- mkPMU(2);
    Operation_IFC mod_122_inner = mod_122_bufferize.operation;
    Operation_IFC mod_122 <- mkDebugOperation(mod_122_inner, "mod_122");
    rule rule_107;
        ChannelMessage t;
        t <- mod_83.get(0);
        mod_84.put(0, t);
    endrule
    rule rule_108;
        ChannelMessage t;
        t <- mod_122.get(1);
        mod_86.put(1, t);
    endrule
    rule rule_109;
        ChannelMessage t;
        t <- mod_117.get(0);
        mod_116.put(1, t);
    endrule
    rule rule_110;
        ChannelMessage t;
        t <- mod_115.get(0);
        mod_114.put(1, t);
    endrule
    rule rule_111;
        ChannelMessage t;
        t <- mod_85.get(0);
        mod_86.put(0, t);
    endrule
    rule rule_112;
        ChannelMessage t;
        t <- mod_90.get(0);
        mod_120.put(0, t);
    endrule
    rule rule_113;
        ChannelMessage t;
        t <- mod_100.get(1);
        mod_98.put(1, t);
    endrule
    rule rule_114;
        ChannelMessage t;
        t <- mod_110.get(0);
        mod_111.put(0, t);
    endrule
    rule rule_115;
        ChannelMessage t;
        t <- mod_101.get(1);
        mod_97.put(1, t);
    endrule
    rule rule_116;
        ChannelMessage t;
        t <- mod_107.get(0);
        mod_93.put(1, t);
    endrule
    rule rule_117;
        ChannelMessage t;
        t <- mod_105.get(0);
        mod_104.put(0, t);
    endrule
    rule rule_118;
        ChannelMessage t;
        t <- mod_98.get(1);
        mod_99.put(1, t);
    endrule
    rule rule_119;
        ChannelMessage t;
        t <- mod_116.get(1);
        mod_91.put(1, t);
    endrule
    rule rule_120;
        ChannelMessage t;
        t <- mod_94.get(1);
        mod_95.put(0, t);
    endrule
    rule rule_121;
        ChannelMessage t;
        t <- mod_92.get(0);
        mod_93.put(0, t);
    endrule
    rule rule_122;
        ChannelMessage t;
        t <- mod_102.get(1);
        mod_95.put(1, t);
    endrule
    rule rule_123;
        ChannelMessage t;
        t <- mod_89.get(0);
        mod_114.put(0, t);
    endrule
    rule rule_124;
        ChannelMessage t;
        t <- mod_114.get(1);
        mod_109.put(0, t);
    endrule
    rule rule_125;
        ChannelMessage t;
        t <- mod_119.get(0);
        mod_118.put(0, t);
    endrule
    rule rule_126;
        ChannelMessage t;
        t <- mod_102.get(0);
        mod_103.put(0, t);
    endrule
    rule rule_127;
        ChannelMessage t;
        t <- mod_84.get(0);
        mod_85.put(0, t);
    endrule
    rule rule_128;
        ChannelMessage t;
        t <- mod_95.get(0);
        mod_96.put(0, t);
    endrule
    rule rule_129;
        ChannelMessage t;
        t <- mod_101.get(0);
        mod_101.put(1, t);
    endrule
    rule rule_130;
        ChannelMessage t;
        t <- mod_120.get(0);
        mod_90.put(1, t);
    endrule
    rule rule_131;
        ChannelMessage t;
        t <- mod_86.get(0);
        mod_122.put(0, t);
    endrule
    rule rule_132;
        ChannelMessage t;
        t <- mod_104.get(0);
        mod_102.put(0, t);
    endrule
    rule rule_133;
        ChannelMessage t;
        t <- mod_96.get(0);
        mod_97.put(0, t);
    endrule
    rule rule_134;
        ChannelMessage t;
        t <- mod_91.get(0);
        mod_92.put(0, t);
    endrule
    rule rule_135;
        ChannelMessage t;
        t <- mod_116.get(0);
        mod_117.put(0, t);
    endrule
    rule rule_136;
        ChannelMessage t;
        t <- mod_111.get(0);
        mod_110.put(1, t);
    endrule
    rule rule_137;
        ChannelMessage t;
        t <- mod_113.get(0);
        mod_112.put(0, t);
    endrule
    rule rule_138;
        ChannelMessage t;
        t <- mod_88.get(0);
        mod_121.put(0, t);
    endrule
    rule rule_139;
        ChannelMessage t;
        t <- mod_87.get(3);
        mod_88.put(0, t);
    endrule
    rule rule_140;
        ChannelMessage t;
        t <- mod_100.get(0);
        mod_100.put(1, t);
    endrule
    rule rule_141;
        ChannelMessage t;
        t <- mod_108.get(0);
        mod_107.put(0, t);
    endrule
    rule rule_142;
        ChannelMessage t;
        t <- mod_88.get(1);
        mod_89.put(0, t);
    endrule
    rule rule_143;
        ChannelMessage t;
        t <- mod_97.get(0);
        mod_101.put(0, t);
    endrule
    rule rule_144;
        ChannelMessage t;
        t <- mod_86.get(1);
        mod_87.put(0, t);
    endrule
    rule rule_145;
        ChannelMessage t;
        t <- mod_106.get(0);
        mod_94.put(1, t);
    endrule
    rule rule_146;
        ChannelMessage t;
        t <- mod_109.get(0);
        mod_108.put(0, t);
    endrule
    rule rule_147;
        ChannelMessage t;
        t <- mod_94.get(0);
        mod_106.put(0, t);
    endrule
    rule rule_148;
        ChannelMessage t;
        t <- mod_114.get(0);
        mod_115.put(0, t);
    endrule
    rule rule_149;
        ChannelMessage t;
        t <- mod_90.get(1);
        mod_91.put(0, t);
    endrule
    rule rule_150;
        ChannelMessage t;
        t <- mod_93.get(0);
        mod_94.put(0, t);
    endrule
    rule rule_151;
        ChannelMessage t;
        t <- mod_121.get(0);
        mod_88.put(1, t);
    endrule
    rule rule_152;
        ChannelMessage t;
        t <- mod_98.get(0);
        mod_100.put(0, t);
    endrule
    rule rule_153;
        ChannelMessage t;
        t <- mod_97.get(1);
        mod_98.put(0, t);
    endrule
    rule rule_154;
        ChannelMessage t;
        t <- mod_103.get(0);
        mod_102.put(1, t);
    endrule
    rule rule_155;
        ChannelMessage t;
        t <- mod_89.get(1);
        mod_90.put(0, t);
    endrule
    rule rule_156;
        ChannelMessage t;
        t <- mod_110.get(1);
        mod_109.put(1, t);
    endrule
    rule rule_157;
        ChannelMessage t;
        t <- mod_118.get(0);
        mod_116.put(0, t);
    endrule
    rule rule_158;
        ChannelMessage t;
        t <- mod_112.get(0);
        mod_110.put(0, t);
    endrule
    rule rule_159;
        ChannelMessage t;
        t <- mod_122.get(0);
        mod_122.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_83.put(0, t);
        end
        if (i == 1) begin
            mod_99.put(0, t);
        end
        if (i == 2) begin
            mod_105.put(0, t);
        end
        if (i == 3) begin
            mod_113.put(0, t);
        end
        if (i == 4) begin
            mod_119.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_87.get(0);
        end
        if (i == 0) begin
            t <- mod_87.get(1);
        end
        if (i == 3) begin
            t <- mod_87.get(2);
        end
        if (i == 2) begin
            t <- mod_99.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6037 (Operation_IFC);
    Operation_IFC mod_124_inner <- mkReshape(2, 64);
    Operation_IFC mod_124 <- mkDebugOperation(mod_124_inner, "mod_124");
    Operation_IFC mod_125_inner <- mkFlatten(1);
    Operation_IFC mod_125 <- mkDebugOperation(mod_125_inner, "mod_125");
    Operation_IFC mod_126_inner <- mkFlatten(2);
    Operation_IFC mod_126 <- mkDebugOperation(mod_126_inner, "mod_126");
    Operation_IFC mod_127_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_127 <- mkDebugOperation(mod_127_inner, "mod_127");
    Broadcast_IFC#(4) mod_128_inner <- mkBroadcast(4);
    Operation_IFC mod_128 <- mkDebugOperation(mod_128_inner.op, "mod_128");
    PMU_IFC mod_129_bufferize <- mkPMU(2);
    Operation_IFC mod_129_inner = mod_129_bufferize.operation;
    Operation_IFC mod_129 <- mkDebugOperation(mod_129_inner, "mod_129");
    Broadcast_IFC#(2) mod_130_inner <- mkBroadcast(2);
    Operation_IFC mod_130 <- mkDebugOperation(mod_130_inner.op, "mod_130");
    PMU_IFC mod_131_bufferize <- mkPMU(1);
    Operation_IFC mod_131_inner = mod_131_bufferize.operation;
    Operation_IFC mod_131 <- mkDebugOperation(mod_131_inner, "mod_131");
    Operation_IFC mod_132_inner <- mkBinaryMap(1153, matmul_t_tile);
    Operation_IFC mod_132 <- mkDebugOperation(mod_132_inner, "mod_132");
    Operation_IFC mod_133_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_133 <- mkDebugOperation(mod_133_inner, "mod_133");
    Operation_IFC mod_134_inner <- mkBinaryMap(1921, mul_tile);
    Operation_IFC mod_134 <- mkDebugOperation(mod_134_inner, "mod_134");
    PMU_IFC mod_135_bufferize <- mkPMU(1);
    Operation_IFC mod_135_inner = mod_135_bufferize.operation;
    Operation_IFC mod_135 <- mkDebugOperation(mod_135_inner, "mod_135");
    Operation_IFC mod_136_inner <- mkBinaryMap(2557, matmul_t_tile);
    Operation_IFC mod_136 <- mkDebugOperation(mod_136_inner, "mod_136");
    Operation_IFC mod_137_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_137 <- mkDebugOperation(mod_137_inner, "mod_137");
    Operation_IFC mod_138_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_138 <- mkDebugOperation(mod_138_inner, "mod_138");
    Operation_IFC mod_139_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_139 <- mkDebugOperation(mod_139_inner, "mod_139");
    Operation_IFC mod_140_inner <- mkBinaryMap(2820, mul_tile);
    Operation_IFC mod_140 <- mkDebugOperation(mod_140_inner, "mod_140");
    PMU_IFC mod_141_bufferize <- mkPMU(1);
    Operation_IFC mod_141_inner = mod_141_bufferize.operation;
    Operation_IFC mod_141 <- mkDebugOperation(mod_141_inner, "mod_141");
    PMU_IFC mod_142_bufferize <- mkPMU(2);
    Operation_IFC mod_142_inner = mod_142_bufferize.operation;
    Operation_IFC mod_142 <- mkDebugOperation(mod_142_inner, "mod_142");
    PMU_IFC mod_143_bufferize <- mkPMU(2);
    Operation_IFC mod_143_inner = mod_143_bufferize.operation;
    Operation_IFC mod_143 <- mkDebugOperation(mod_143_inner, "mod_143");
    Operation_IFC mod_144_inner <- mkRepeatStatic(8);
    Operation_IFC mod_144 <- mkDebugOperation(mod_144_inner, "mod_144");
    Operation_IFC mod_145_inner <- mkFlatten(1);
    Operation_IFC mod_145 <- mkDebugOperation(mod_145_inner, "mod_145");
    Operation_IFC mod_146_inner <- mkFlatten(0);
    Operation_IFC mod_146 <- mkDebugOperation(mod_146_inner, "mod_146");
    Operation_IFC mod_147_inner <- mkRepeatStatic(3);
    Operation_IFC mod_147 <- mkDebugOperation(mod_147_inner, "mod_147");
    Operation_IFC mod_148_inner <- mkUnaryMap(1793, silu_tile);
    Operation_IFC mod_148 <- mkDebugOperation(mod_148_inner, "mod_148");
    Operation_IFC mod_149_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_149 <- mkDebugOperation(mod_149_inner, "mod_149");
    Operation_IFC mod_150_inner <- mkBinaryMap(1665, matmul_t_tile);
    Operation_IFC mod_150 <- mkDebugOperation(mod_150_inner, "mod_150");
    PMU_IFC mod_151_bufferize <- mkPMU(2);
    Operation_IFC mod_151_inner = mod_151_bufferize.operation;
    Operation_IFC mod_151 <- mkDebugOperation(mod_151_inner, "mod_151");
    Operation_IFC mod_152_inner <- mkRepeatStatic(8);
    Operation_IFC mod_152 <- mkDebugOperation(mod_152_inner, "mod_152");
    Operation_IFC mod_153_inner <- mkFlatten(1);
    Operation_IFC mod_153 <- mkDebugOperation(mod_153_inner, "mod_153");
    Operation_IFC mod_154_inner <- mkFlatten(0);
    Operation_IFC mod_154 <- mkDebugOperation(mod_154_inner, "mod_154");
    PMU_IFC mod_155_bufferize <- mkPMU(1);
    Operation_IFC mod_155_inner = mod_155_bufferize.operation;
    Operation_IFC mod_155 <- mkDebugOperation(mod_155_inner, "mod_155");
    Operation_IFC mod_156_inner <- mkRepeatStatic(16);
    Operation_IFC mod_156 <- mkDebugOperation(mod_156_inner, "mod_156");
    PMU_IFC mod_157_bufferize <- mkPMU(2);
    Operation_IFC mod_157_inner = mod_157_bufferize.operation;
    Operation_IFC mod_157 <- mkDebugOperation(mod_157_inner, "mod_157");
    Operation_IFC mod_158_inner <- mkRepeatStatic(8);
    Operation_IFC mod_158 <- mkDebugOperation(mod_158_inner, "mod_158");
    Operation_IFC mod_159_inner <- mkFlatten(1);
    Operation_IFC mod_159 <- mkDebugOperation(mod_159_inner, "mod_159");
    Operation_IFC mod_160_inner <- mkFlatten(0);
    Operation_IFC mod_160 <- mkDebugOperation(mod_160_inner, "mod_160");
    Operation_IFC mod_161_inner <- mkRepeatStatic(16);
    Operation_IFC mod_161 <- mkDebugOperation(mod_161_inner, "mod_161");
    Operation_IFC mod_162_inner <- mkRepeatStatic(2);
    Operation_IFC mod_162 <- mkDebugOperation(mod_162_inner, "mod_162");
    PMU_IFC mod_163_bufferize <- mkPMU(2);
    Operation_IFC mod_163_inner = mod_163_bufferize.operation;
    Operation_IFC mod_163 <- mkDebugOperation(mod_163_inner, "mod_163");
    rule rule_160;
        ChannelMessage t;
        t <- mod_135.get(1);
        mod_136.put(0, t);
    endrule
    rule rule_161;
        ChannelMessage t;
        t <- mod_139.get(1);
        mod_140.put(1, t);
    endrule
    rule rule_162;
        ChannelMessage t;
        t <- mod_141.get(1);
        mod_139.put(1, t);
    endrule
    rule rule_163;
        ChannelMessage t;
        t <- mod_132.get(0);
        mod_133.put(0, t);
    endrule
    rule rule_164;
        ChannelMessage t;
        t <- mod_136.get(0);
        mod_137.put(0, t);
    endrule
    rule rule_165;
        ChannelMessage t;
        t <- mod_141.get(0);
        mod_141.put(1, t);
    endrule
    rule rule_166;
        ChannelMessage t;
        t <- mod_143.get(1);
        mod_136.put(1, t);
    endrule
    rule rule_167;
        ChannelMessage t;
        t <- mod_147.get(0);
        mod_135.put(1, t);
    endrule
    rule rule_168;
        ChannelMessage t;
        t <- mod_157.get(1);
        mod_132.put(1, t);
    endrule
    rule rule_169;
        ChannelMessage t;
        t <- mod_131.get(1);
        mod_132.put(0, t);
    endrule
    rule rule_170;
        ChannelMessage t;
        t <- mod_139.get(0);
        mod_141.put(0, t);
    endrule
    rule rule_171;
        ChannelMessage t;
        t <- mod_138.get(0);
        mod_142.put(0, t);
    endrule
    rule rule_172;
        ChannelMessage t;
        t <- mod_163.get(1);
        mod_127.put(1, t);
    endrule
    rule rule_173;
        ChannelMessage t;
        t <- mod_152.get(0);
        mod_151.put(1, t);
    endrule
    rule rule_174;
        ChannelMessage t;
        t <- mod_135.get(0);
        mod_147.put(0, t);
    endrule
    rule rule_175;
        ChannelMessage t;
        t <- mod_127.get(1);
        mod_128.put(0, t);
    endrule
    rule rule_176;
        ChannelMessage t;
        t <- mod_128.get(3);
        mod_129.put(0, t);
    endrule
    rule rule_177;
        ChannelMessage t;
        t <- mod_146.get(0);
        mod_145.put(0, t);
    endrule
    rule rule_178;
        ChannelMessage t;
        t <- mod_151.get(0);
        mod_152.put(0, t);
    endrule
    rule rule_179;
        ChannelMessage t;
        t <- mod_155.get(0);
        mod_156.put(0, t);
    endrule
    rule rule_180;
        ChannelMessage t;
        t <- mod_134.get(0);
        mod_135.put(0, t);
    endrule
    rule rule_181;
        ChannelMessage t;
        t <- mod_126.get(0);
        mod_127.put(0, t);
    endrule
    rule rule_182;
        ChannelMessage t;
        t <- mod_129.get(1);
        mod_130.put(0, t);
    endrule
    rule rule_183;
        ChannelMessage t;
        t <- mod_130.get(1);
        mod_131.put(0, t);
    endrule
    rule rule_184;
        ChannelMessage t;
        t <- mod_144.get(0);
        mod_143.put(1, t);
    endrule
    rule rule_185;
        ChannelMessage t;
        t <- mod_154.get(0);
        mod_153.put(0, t);
    endrule
    rule rule_186;
        ChannelMessage t;
        t <- mod_137.get(0);
        mod_138.put(0, t);
    endrule
    rule rule_187;
        ChannelMessage t;
        t <- mod_131.get(0);
        mod_161.put(0, t);
    endrule
    rule rule_188;
        ChannelMessage t;
        t <- mod_138.get(1);
        mod_139.put(0, t);
    endrule
    rule rule_189;
        ChannelMessage t;
        t <- mod_127.get(0);
        mod_163.put(0, t);
    endrule
    rule rule_190;
        ChannelMessage t;
        t <- mod_142.get(0);
        mod_142.put(1, t);
    endrule
    rule rule_191;
        ChannelMessage t;
        t <- mod_145.get(0);
        mod_143.put(0, t);
    endrule
    rule rule_192;
        ChannelMessage t;
        t <- mod_160.get(0);
        mod_159.put(0, t);
    endrule
    rule rule_193;
        ChannelMessage t;
        t <- mod_155.get(1);
        mod_150.put(0, t);
    endrule
    rule rule_194;
        ChannelMessage t;
        t <- mod_133.get(0);
        mod_134.put(0, t);
    endrule
    rule rule_195;
        ChannelMessage t;
        t <- mod_149.get(0);
        mod_148.put(0, t);
    endrule
    rule rule_196;
        ChannelMessage t;
        t <- mod_124.get(0);
        mod_125.put(0, t);
    endrule
    rule rule_197;
        ChannelMessage t;
        t <- mod_142.get(1);
        mod_138.put(1, t);
    endrule
    rule rule_198;
        ChannelMessage t;
        t <- mod_130.get(0);
        mod_155.put(0, t);
    endrule
    rule rule_199;
        ChannelMessage t;
        t <- mod_159.get(0);
        mod_157.put(0, t);
    endrule
    rule rule_200;
        ChannelMessage t;
        t <- mod_162.get(0);
        mod_129.put(1, t);
    endrule
    rule rule_201;
        ChannelMessage t;
        t <- mod_157.get(0);
        mod_158.put(0, t);
    endrule
    rule rule_202;
        ChannelMessage t;
        t <- mod_151.get(1);
        mod_150.put(1, t);
    endrule
    rule rule_203;
        ChannelMessage t;
        t <- mod_156.get(0);
        mod_155.put(1, t);
    endrule
    rule rule_204;
        ChannelMessage t;
        t <- mod_163.get(0);
        mod_163.put(1, t);
    endrule
    rule rule_205;
        ChannelMessage t;
        t <- mod_150.get(0);
        mod_149.put(0, t);
    endrule
    rule rule_206;
        ChannelMessage t;
        t <- mod_158.get(0);
        mod_157.put(1, t);
    endrule
    rule rule_207;
        ChannelMessage t;
        t <- mod_153.get(0);
        mod_151.put(0, t);
    endrule
    rule rule_208;
        ChannelMessage t;
        t <- mod_143.get(0);
        mod_144.put(0, t);
    endrule
    rule rule_209;
        ChannelMessage t;
        t <- mod_148.get(0);
        mod_134.put(1, t);
    endrule
    rule rule_210;
        ChannelMessage t;
        t <- mod_125.get(0);
        mod_126.put(0, t);
    endrule
    rule rule_211;
        ChannelMessage t;
        t <- mod_161.get(0);
        mod_131.put(1, t);
    endrule
    rule rule_212;
        ChannelMessage t;
        t <- mod_129.get(0);
        mod_162.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_124.put(0, t);
        end
        if (i == 1) begin
            mod_140.put(0, t);
        end
        if (i == 2) begin
            mod_146.put(0, t);
        end
        if (i == 3) begin
            mod_154.put(0, t);
        end
        if (i == 4) begin
            mod_160.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_128.get(0);
        end
        if (i == 2) begin
            t <- mod_128.get(1);
        end
        if (i == 1) begin
            t <- mod_128.get(2);
        end
        if (i == 0) begin
            t <- mod_140.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6038 (Operation_IFC);
    Operation_IFC mod_165_inner <- mkReshape(2, 64);
    Operation_IFC mod_165 <- mkDebugOperation(mod_165_inner, "mod_165");
    Operation_IFC mod_166_inner <- mkFlatten(1);
    Operation_IFC mod_166 <- mkDebugOperation(mod_166_inner, "mod_166");
    Operation_IFC mod_167_inner <- mkFlatten(2);
    Operation_IFC mod_167 <- mkDebugOperation(mod_167_inner, "mod_167");
    Operation_IFC mod_168_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_168 <- mkDebugOperation(mod_168_inner, "mod_168");
    Broadcast_IFC#(4) mod_169_inner <- mkBroadcast(4);
    Operation_IFC mod_169 <- mkDebugOperation(mod_169_inner.op, "mod_169");
    PMU_IFC mod_170_bufferize <- mkPMU(2);
    Operation_IFC mod_170_inner = mod_170_bufferize.operation;
    Operation_IFC mod_170 <- mkDebugOperation(mod_170_inner, "mod_170");
    Broadcast_IFC#(2) mod_171_inner <- mkBroadcast(2);
    Operation_IFC mod_171 <- mkDebugOperation(mod_171_inner.op, "mod_171");
    PMU_IFC mod_172_bufferize <- mkPMU(1);
    Operation_IFC mod_172_inner = mod_172_bufferize.operation;
    Operation_IFC mod_172 <- mkDebugOperation(mod_172_inner, "mod_172");
    Operation_IFC mod_173_inner <- mkBinaryMap(1152, matmul_t_tile);
    Operation_IFC mod_173 <- mkDebugOperation(mod_173_inner, "mod_173");
    Operation_IFC mod_174_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_174 <- mkDebugOperation(mod_174_inner, "mod_174");
    Operation_IFC mod_175_inner <- mkBinaryMap(1920, mul_tile);
    Operation_IFC mod_175 <- mkDebugOperation(mod_175_inner, "mod_175");
    PMU_IFC mod_176_bufferize <- mkPMU(1);
    Operation_IFC mod_176_inner = mod_176_bufferize.operation;
    Operation_IFC mod_176 <- mkDebugOperation(mod_176_inner, "mod_176");
    Operation_IFC mod_177_inner <- mkBinaryMap(2555, matmul_t_tile);
    Operation_IFC mod_177 <- mkDebugOperation(mod_177_inner, "mod_177");
    Operation_IFC mod_178_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_178 <- mkDebugOperation(mod_178_inner, "mod_178");
    Operation_IFC mod_179_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_179 <- mkDebugOperation(mod_179_inner, "mod_179");
    Operation_IFC mod_180_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_180 <- mkDebugOperation(mod_180_inner, "mod_180");
    Operation_IFC mod_181_inner <- mkBinaryMap(2819, mul_tile);
    Operation_IFC mod_181 <- mkDebugOperation(mod_181_inner, "mod_181");
    PMU_IFC mod_182_bufferize <- mkPMU(1);
    Operation_IFC mod_182_inner = mod_182_bufferize.operation;
    Operation_IFC mod_182 <- mkDebugOperation(mod_182_inner, "mod_182");
    PMU_IFC mod_183_bufferize <- mkPMU(2);
    Operation_IFC mod_183_inner = mod_183_bufferize.operation;
    Operation_IFC mod_183 <- mkDebugOperation(mod_183_inner, "mod_183");
    PMU_IFC mod_184_bufferize <- mkPMU(2);
    Operation_IFC mod_184_inner = mod_184_bufferize.operation;
    Operation_IFC mod_184 <- mkDebugOperation(mod_184_inner, "mod_184");
    Operation_IFC mod_185_inner <- mkRepeatStatic(8);
    Operation_IFC mod_185 <- mkDebugOperation(mod_185_inner, "mod_185");
    Operation_IFC mod_186_inner <- mkFlatten(1);
    Operation_IFC mod_186 <- mkDebugOperation(mod_186_inner, "mod_186");
    Operation_IFC mod_187_inner <- mkFlatten(0);
    Operation_IFC mod_187 <- mkDebugOperation(mod_187_inner, "mod_187");
    Operation_IFC mod_188_inner <- mkRepeatStatic(3);
    Operation_IFC mod_188 <- mkDebugOperation(mod_188_inner, "mod_188");
    Operation_IFC mod_189_inner <- mkUnaryMap(1792, silu_tile);
    Operation_IFC mod_189 <- mkDebugOperation(mod_189_inner, "mod_189");
    Operation_IFC mod_190_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_190 <- mkDebugOperation(mod_190_inner, "mod_190");
    Operation_IFC mod_191_inner <- mkBinaryMap(1664, matmul_t_tile);
    Operation_IFC mod_191 <- mkDebugOperation(mod_191_inner, "mod_191");
    PMU_IFC mod_192_bufferize <- mkPMU(2);
    Operation_IFC mod_192_inner = mod_192_bufferize.operation;
    Operation_IFC mod_192 <- mkDebugOperation(mod_192_inner, "mod_192");
    Operation_IFC mod_193_inner <- mkRepeatStatic(8);
    Operation_IFC mod_193 <- mkDebugOperation(mod_193_inner, "mod_193");
    Operation_IFC mod_194_inner <- mkFlatten(1);
    Operation_IFC mod_194 <- mkDebugOperation(mod_194_inner, "mod_194");
    Operation_IFC mod_195_inner <- mkFlatten(0);
    Operation_IFC mod_195 <- mkDebugOperation(mod_195_inner, "mod_195");
    PMU_IFC mod_196_bufferize <- mkPMU(1);
    Operation_IFC mod_196_inner = mod_196_bufferize.operation;
    Operation_IFC mod_196 <- mkDebugOperation(mod_196_inner, "mod_196");
    Operation_IFC mod_197_inner <- mkRepeatStatic(16);
    Operation_IFC mod_197 <- mkDebugOperation(mod_197_inner, "mod_197");
    PMU_IFC mod_198_bufferize <- mkPMU(2);
    Operation_IFC mod_198_inner = mod_198_bufferize.operation;
    Operation_IFC mod_198 <- mkDebugOperation(mod_198_inner, "mod_198");
    Operation_IFC mod_199_inner <- mkRepeatStatic(8);
    Operation_IFC mod_199 <- mkDebugOperation(mod_199_inner, "mod_199");
    Operation_IFC mod_200_inner <- mkFlatten(1);
    Operation_IFC mod_200 <- mkDebugOperation(mod_200_inner, "mod_200");
    Operation_IFC mod_201_inner <- mkFlatten(0);
    Operation_IFC mod_201 <- mkDebugOperation(mod_201_inner, "mod_201");
    Operation_IFC mod_202_inner <- mkRepeatStatic(16);
    Operation_IFC mod_202 <- mkDebugOperation(mod_202_inner, "mod_202");
    Operation_IFC mod_203_inner <- mkRepeatStatic(2);
    Operation_IFC mod_203 <- mkDebugOperation(mod_203_inner, "mod_203");
    PMU_IFC mod_204_bufferize <- mkPMU(2);
    Operation_IFC mod_204_inner = mod_204_bufferize.operation;
    Operation_IFC mod_204 <- mkDebugOperation(mod_204_inner, "mod_204");
    rule rule_213;
        ChannelMessage t;
        t <- mod_170.get(1);
        mod_171.put(0, t);
    endrule
    rule rule_214;
        ChannelMessage t;
        t <- mod_201.get(0);
        mod_200.put(0, t);
    endrule
    rule rule_215;
        ChannelMessage t;
        t <- mod_184.get(1);
        mod_177.put(1, t);
    endrule
    rule rule_216;
        ChannelMessage t;
        t <- mod_196.get(0);
        mod_197.put(0, t);
    endrule
    rule rule_217;
        ChannelMessage t;
        t <- mod_183.get(1);
        mod_179.put(1, t);
    endrule
    rule rule_218;
        ChannelMessage t;
        t <- mod_187.get(0);
        mod_186.put(0, t);
    endrule
    rule rule_219;
        ChannelMessage t;
        t <- mod_195.get(0);
        mod_194.put(0, t);
    endrule
    rule rule_220;
        ChannelMessage t;
        t <- mod_193.get(0);
        mod_192.put(1, t);
    endrule
    rule rule_221;
        ChannelMessage t;
        t <- mod_188.get(0);
        mod_176.put(1, t);
    endrule
    rule rule_222;
        ChannelMessage t;
        t <- mod_204.get(0);
        mod_204.put(1, t);
    endrule
    rule rule_223;
        ChannelMessage t;
        t <- mod_196.get(1);
        mod_191.put(0, t);
    endrule
    rule rule_224;
        ChannelMessage t;
        t <- mod_199.get(0);
        mod_198.put(1, t);
    endrule
    rule rule_225;
        ChannelMessage t;
        t <- mod_172.get(0);
        mod_202.put(0, t);
    endrule
    rule rule_226;
        ChannelMessage t;
        t <- mod_166.get(0);
        mod_167.put(0, t);
    endrule
    rule rule_227;
        ChannelMessage t;
        t <- mod_173.get(0);
        mod_174.put(0, t);
    endrule
    rule rule_228;
        ChannelMessage t;
        t <- mod_191.get(0);
        mod_190.put(0, t);
    endrule
    rule rule_229;
        ChannelMessage t;
        t <- mod_203.get(0);
        mod_170.put(1, t);
    endrule
    rule rule_230;
        ChannelMessage t;
        t <- mod_182.get(0);
        mod_182.put(1, t);
    endrule
    rule rule_231;
        ChannelMessage t;
        t <- mod_186.get(0);
        mod_184.put(0, t);
    endrule
    rule rule_232;
        ChannelMessage t;
        t <- mod_180.get(0);
        mod_182.put(0, t);
    endrule
    rule rule_233;
        ChannelMessage t;
        t <- mod_167.get(0);
        mod_168.put(0, t);
    endrule
    rule rule_234;
        ChannelMessage t;
        t <- mod_200.get(0);
        mod_198.put(0, t);
    endrule
    rule rule_235;
        ChannelMessage t;
        t <- mod_197.get(0);
        mod_196.put(1, t);
    endrule
    rule rule_236;
        ChannelMessage t;
        t <- mod_176.get(1);
        mod_177.put(0, t);
    endrule
    rule rule_237;
        ChannelMessage t;
        t <- mod_179.get(1);
        mod_180.put(0, t);
    endrule
    rule rule_238;
        ChannelMessage t;
        t <- mod_177.get(0);
        mod_178.put(0, t);
    endrule
    rule rule_239;
        ChannelMessage t;
        t <- mod_185.get(0);
        mod_184.put(1, t);
    endrule
    rule rule_240;
        ChannelMessage t;
        t <- mod_198.get(1);
        mod_173.put(1, t);
    endrule
    rule rule_241;
        ChannelMessage t;
        t <- mod_192.get(0);
        mod_193.put(0, t);
    endrule
    rule rule_242;
        ChannelMessage t;
        t <- mod_184.get(0);
        mod_185.put(0, t);
    endrule
    rule rule_243;
        ChannelMessage t;
        t <- mod_194.get(0);
        mod_192.put(0, t);
    endrule
    rule rule_244;
        ChannelMessage t;
        t <- mod_179.get(0);
        mod_183.put(0, t);
    endrule
    rule rule_245;
        ChannelMessage t;
        t <- mod_183.get(0);
        mod_183.put(1, t);
    endrule
    rule rule_246;
        ChannelMessage t;
        t <- mod_182.get(1);
        mod_180.put(1, t);
    endrule
    rule rule_247;
        ChannelMessage t;
        t <- mod_172.get(1);
        mod_173.put(0, t);
    endrule
    rule rule_248;
        ChannelMessage t;
        t <- mod_189.get(0);
        mod_175.put(1, t);
    endrule
    rule rule_249;
        ChannelMessage t;
        t <- mod_192.get(1);
        mod_191.put(1, t);
    endrule
    rule rule_250;
        ChannelMessage t;
        t <- mod_198.get(0);
        mod_199.put(0, t);
    endrule
    rule rule_251;
        ChannelMessage t;
        t <- mod_165.get(0);
        mod_166.put(0, t);
    endrule
    rule rule_252;
        ChannelMessage t;
        t <- mod_168.get(1);
        mod_169.put(0, t);
    endrule
    rule rule_253;
        ChannelMessage t;
        t <- mod_202.get(0);
        mod_172.put(1, t);
    endrule
    rule rule_254;
        ChannelMessage t;
        t <- mod_204.get(1);
        mod_168.put(1, t);
    endrule
    rule rule_255;
        ChannelMessage t;
        t <- mod_171.get(1);
        mod_172.put(0, t);
    endrule
    rule rule_256;
        ChannelMessage t;
        t <- mod_176.get(0);
        mod_188.put(0, t);
    endrule
    rule rule_257;
        ChannelMessage t;
        t <- mod_178.get(0);
        mod_179.put(0, t);
    endrule
    rule rule_258;
        ChannelMessage t;
        t <- mod_175.get(0);
        mod_176.put(0, t);
    endrule
    rule rule_259;
        ChannelMessage t;
        t <- mod_168.get(0);
        mod_204.put(0, t);
    endrule
    rule rule_260;
        ChannelMessage t;
        t <- mod_169.get(3);
        mod_170.put(0, t);
    endrule
    rule rule_261;
        ChannelMessage t;
        t <- mod_171.get(0);
        mod_196.put(0, t);
    endrule
    rule rule_262;
        ChannelMessage t;
        t <- mod_180.get(1);
        mod_181.put(1, t);
    endrule
    rule rule_263;
        ChannelMessage t;
        t <- mod_170.get(0);
        mod_203.put(0, t);
    endrule
    rule rule_264;
        ChannelMessage t;
        t <- mod_190.get(0);
        mod_189.put(0, t);
    endrule
    rule rule_265;
        ChannelMessage t;
        t <- mod_174.get(0);
        mod_175.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_165.put(0, t);
        end
        if (i == 1) begin
            mod_181.put(0, t);
        end
        if (i == 2) begin
            mod_187.put(0, t);
        end
        if (i == 3) begin
            mod_195.put(0, t);
        end
        if (i == 4) begin
            mod_201.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_169.get(0);
        end
        if (i == 2) begin
            t <- mod_169.get(1);
        end
        if (i == 0) begin
            t <- mod_169.get(2);
        end
        if (i == 1) begin
            t <- mod_181.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6039 (Operation_IFC);
    Operation_IFC mod_206_inner <- mkReshape(2, 64);
    Operation_IFC mod_206 <- mkDebugOperation(mod_206_inner, "mod_206");
    Operation_IFC mod_207_inner <- mkFlatten(1);
    Operation_IFC mod_207 <- mkDebugOperation(mod_207_inner, "mod_207");
    Operation_IFC mod_208_inner <- mkFlatten(2);
    Operation_IFC mod_208 <- mkDebugOperation(mod_208_inner, "mod_208");
    Operation_IFC mod_209_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_209 <- mkDebugOperation(mod_209_inner, "mod_209");
    Broadcast_IFC#(4) mod_210_inner <- mkBroadcast(4);
    Operation_IFC mod_210 <- mkDebugOperation(mod_210_inner.op, "mod_210");
    PMU_IFC mod_211_bufferize <- mkPMU(2);
    Operation_IFC mod_211_inner = mod_211_bufferize.operation;
    Operation_IFC mod_211 <- mkDebugOperation(mod_211_inner, "mod_211");
    Broadcast_IFC#(2) mod_212_inner <- mkBroadcast(2);
    Operation_IFC mod_212 <- mkDebugOperation(mod_212_inner.op, "mod_212");
    PMU_IFC mod_213_bufferize <- mkPMU(1);
    Operation_IFC mod_213_inner = mod_213_bufferize.operation;
    Operation_IFC mod_213 <- mkDebugOperation(mod_213_inner, "mod_213");
    Operation_IFC mod_214_inner <- mkBinaryMap(1151, matmul_t_tile);
    Operation_IFC mod_214 <- mkDebugOperation(mod_214_inner, "mod_214");
    Operation_IFC mod_215_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_215 <- mkDebugOperation(mod_215_inner, "mod_215");
    Operation_IFC mod_216_inner <- mkBinaryMap(1919, mul_tile);
    Operation_IFC mod_216 <- mkDebugOperation(mod_216_inner, "mod_216");
    PMU_IFC mod_217_bufferize <- mkPMU(1);
    Operation_IFC mod_217_inner = mod_217_bufferize.operation;
    Operation_IFC mod_217 <- mkDebugOperation(mod_217_inner, "mod_217");
    Operation_IFC mod_218_inner <- mkBinaryMap(2553, matmul_t_tile);
    Operation_IFC mod_218 <- mkDebugOperation(mod_218_inner, "mod_218");
    Operation_IFC mod_219_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_219 <- mkDebugOperation(mod_219_inner, "mod_219");
    Operation_IFC mod_220_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_220 <- mkDebugOperation(mod_220_inner, "mod_220");
    Operation_IFC mod_221_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_221 <- mkDebugOperation(mod_221_inner, "mod_221");
    Operation_IFC mod_222_inner <- mkBinaryMap(2818, mul_tile);
    Operation_IFC mod_222 <- mkDebugOperation(mod_222_inner, "mod_222");
    PMU_IFC mod_223_bufferize <- mkPMU(1);
    Operation_IFC mod_223_inner = mod_223_bufferize.operation;
    Operation_IFC mod_223 <- mkDebugOperation(mod_223_inner, "mod_223");
    PMU_IFC mod_224_bufferize <- mkPMU(2);
    Operation_IFC mod_224_inner = mod_224_bufferize.operation;
    Operation_IFC mod_224 <- mkDebugOperation(mod_224_inner, "mod_224");
    PMU_IFC mod_225_bufferize <- mkPMU(2);
    Operation_IFC mod_225_inner = mod_225_bufferize.operation;
    Operation_IFC mod_225 <- mkDebugOperation(mod_225_inner, "mod_225");
    Operation_IFC mod_226_inner <- mkRepeatStatic(8);
    Operation_IFC mod_226 <- mkDebugOperation(mod_226_inner, "mod_226");
    Operation_IFC mod_227_inner <- mkFlatten(1);
    Operation_IFC mod_227 <- mkDebugOperation(mod_227_inner, "mod_227");
    Operation_IFC mod_228_inner <- mkFlatten(0);
    Operation_IFC mod_228 <- mkDebugOperation(mod_228_inner, "mod_228");
    Operation_IFC mod_229_inner <- mkRepeatStatic(3);
    Operation_IFC mod_229 <- mkDebugOperation(mod_229_inner, "mod_229");
    Operation_IFC mod_230_inner <- mkUnaryMap(1791, silu_tile);
    Operation_IFC mod_230 <- mkDebugOperation(mod_230_inner, "mod_230");
    Operation_IFC mod_231_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_231 <- mkDebugOperation(mod_231_inner, "mod_231");
    Operation_IFC mod_232_inner <- mkBinaryMap(1663, matmul_t_tile);
    Operation_IFC mod_232 <- mkDebugOperation(mod_232_inner, "mod_232");
    PMU_IFC mod_233_bufferize <- mkPMU(2);
    Operation_IFC mod_233_inner = mod_233_bufferize.operation;
    Operation_IFC mod_233 <- mkDebugOperation(mod_233_inner, "mod_233");
    Operation_IFC mod_234_inner <- mkRepeatStatic(8);
    Operation_IFC mod_234 <- mkDebugOperation(mod_234_inner, "mod_234");
    Operation_IFC mod_235_inner <- mkFlatten(1);
    Operation_IFC mod_235 <- mkDebugOperation(mod_235_inner, "mod_235");
    Operation_IFC mod_236_inner <- mkFlatten(0);
    Operation_IFC mod_236 <- mkDebugOperation(mod_236_inner, "mod_236");
    PMU_IFC mod_237_bufferize <- mkPMU(1);
    Operation_IFC mod_237_inner = mod_237_bufferize.operation;
    Operation_IFC mod_237 <- mkDebugOperation(mod_237_inner, "mod_237");
    Operation_IFC mod_238_inner <- mkRepeatStatic(16);
    Operation_IFC mod_238 <- mkDebugOperation(mod_238_inner, "mod_238");
    PMU_IFC mod_239_bufferize <- mkPMU(2);
    Operation_IFC mod_239_inner = mod_239_bufferize.operation;
    Operation_IFC mod_239 <- mkDebugOperation(mod_239_inner, "mod_239");
    Operation_IFC mod_240_inner <- mkRepeatStatic(8);
    Operation_IFC mod_240 <- mkDebugOperation(mod_240_inner, "mod_240");
    Operation_IFC mod_241_inner <- mkFlatten(1);
    Operation_IFC mod_241 <- mkDebugOperation(mod_241_inner, "mod_241");
    Operation_IFC mod_242_inner <- mkFlatten(0);
    Operation_IFC mod_242 <- mkDebugOperation(mod_242_inner, "mod_242");
    Operation_IFC mod_243_inner <- mkRepeatStatic(16);
    Operation_IFC mod_243 <- mkDebugOperation(mod_243_inner, "mod_243");
    Operation_IFC mod_244_inner <- mkRepeatStatic(2);
    Operation_IFC mod_244 <- mkDebugOperation(mod_244_inner, "mod_244");
    PMU_IFC mod_245_bufferize <- mkPMU(2);
    Operation_IFC mod_245_inner = mod_245_bufferize.operation;
    Operation_IFC mod_245 <- mkDebugOperation(mod_245_inner, "mod_245");
    rule rule_266;
        ChannelMessage t;
        t <- mod_239.get(1);
        mod_214.put(1, t);
    endrule
    rule rule_267;
        ChannelMessage t;
        t <- mod_245.get(1);
        mod_209.put(1, t);
    endrule
    rule rule_268;
        ChannelMessage t;
        t <- mod_208.get(0);
        mod_209.put(0, t);
    endrule
    rule rule_269;
        ChannelMessage t;
        t <- mod_218.get(0);
        mod_219.put(0, t);
    endrule
    rule rule_270;
        ChannelMessage t;
        t <- mod_219.get(0);
        mod_220.put(0, t);
    endrule
    rule rule_271;
        ChannelMessage t;
        t <- mod_232.get(0);
        mod_231.put(0, t);
    endrule
    rule rule_272;
        ChannelMessage t;
        t <- mod_226.get(0);
        mod_225.put(1, t);
    endrule
    rule rule_273;
        ChannelMessage t;
        t <- mod_217.get(0);
        mod_229.put(0, t);
    endrule
    rule rule_274;
        ChannelMessage t;
        t <- mod_225.get(0);
        mod_226.put(0, t);
    endrule
    rule rule_275;
        ChannelMessage t;
        t <- mod_244.get(0);
        mod_211.put(1, t);
    endrule
    rule rule_276;
        ChannelMessage t;
        t <- mod_206.get(0);
        mod_207.put(0, t);
    endrule
    rule rule_277;
        ChannelMessage t;
        t <- mod_229.get(0);
        mod_217.put(1, t);
    endrule
    rule rule_278;
        ChannelMessage t;
        t <- mod_241.get(0);
        mod_239.put(0, t);
    endrule
    rule rule_279;
        ChannelMessage t;
        t <- mod_221.get(1);
        mod_222.put(1, t);
    endrule
    rule rule_280;
        ChannelMessage t;
        t <- mod_223.get(1);
        mod_221.put(1, t);
    endrule
    rule rule_281;
        ChannelMessage t;
        t <- mod_224.get(1);
        mod_220.put(1, t);
    endrule
    rule rule_282;
        ChannelMessage t;
        t <- mod_237.get(0);
        mod_238.put(0, t);
    endrule
    rule rule_283;
        ChannelMessage t;
        t <- mod_239.get(0);
        mod_240.put(0, t);
    endrule
    rule rule_284;
        ChannelMessage t;
        t <- mod_211.get(1);
        mod_212.put(0, t);
    endrule
    rule rule_285;
        ChannelMessage t;
        t <- mod_240.get(0);
        mod_239.put(1, t);
    endrule
    rule rule_286;
        ChannelMessage t;
        t <- mod_243.get(0);
        mod_213.put(1, t);
    endrule
    rule rule_287;
        ChannelMessage t;
        t <- mod_209.get(0);
        mod_245.put(0, t);
    endrule
    rule rule_288;
        ChannelMessage t;
        t <- mod_210.get(3);
        mod_211.put(0, t);
    endrule
    rule rule_289;
        ChannelMessage t;
        t <- mod_233.get(0);
        mod_234.put(0, t);
    endrule
    rule rule_290;
        ChannelMessage t;
        t <- mod_213.get(1);
        mod_214.put(0, t);
    endrule
    rule rule_291;
        ChannelMessage t;
        t <- mod_220.get(1);
        mod_221.put(0, t);
    endrule
    rule rule_292;
        ChannelMessage t;
        t <- mod_230.get(0);
        mod_216.put(1, t);
    endrule
    rule rule_293;
        ChannelMessage t;
        t <- mod_225.get(1);
        mod_218.put(1, t);
    endrule
    rule rule_294;
        ChannelMessage t;
        t <- mod_224.get(0);
        mod_224.put(1, t);
    endrule
    rule rule_295;
        ChannelMessage t;
        t <- mod_235.get(0);
        mod_233.put(0, t);
    endrule
    rule rule_296;
        ChannelMessage t;
        t <- mod_237.get(1);
        mod_232.put(0, t);
    endrule
    rule rule_297;
        ChannelMessage t;
        t <- mod_223.get(0);
        mod_223.put(1, t);
    endrule
    rule rule_298;
        ChannelMessage t;
        t <- mod_211.get(0);
        mod_244.put(0, t);
    endrule
    rule rule_299;
        ChannelMessage t;
        t <- mod_233.get(1);
        mod_232.put(1, t);
    endrule
    rule rule_300;
        ChannelMessage t;
        t <- mod_242.get(0);
        mod_241.put(0, t);
    endrule
    rule rule_301;
        ChannelMessage t;
        t <- mod_220.get(0);
        mod_224.put(0, t);
    endrule
    rule rule_302;
        ChannelMessage t;
        t <- mod_212.get(0);
        mod_237.put(0, t);
    endrule
    rule rule_303;
        ChannelMessage t;
        t <- mod_207.get(0);
        mod_208.put(0, t);
    endrule
    rule rule_304;
        ChannelMessage t;
        t <- mod_212.get(1);
        mod_213.put(0, t);
    endrule
    rule rule_305;
        ChannelMessage t;
        t <- mod_214.get(0);
        mod_215.put(0, t);
    endrule
    rule rule_306;
        ChannelMessage t;
        t <- mod_216.get(0);
        mod_217.put(0, t);
    endrule
    rule rule_307;
        ChannelMessage t;
        t <- mod_217.get(1);
        mod_218.put(0, t);
    endrule
    rule rule_308;
        ChannelMessage t;
        t <- mod_227.get(0);
        mod_225.put(0, t);
    endrule
    rule rule_309;
        ChannelMessage t;
        t <- mod_221.get(0);
        mod_223.put(0, t);
    endrule
    rule rule_310;
        ChannelMessage t;
        t <- mod_231.get(0);
        mod_230.put(0, t);
    endrule
    rule rule_311;
        ChannelMessage t;
        t <- mod_238.get(0);
        mod_237.put(1, t);
    endrule
    rule rule_312;
        ChannelMessage t;
        t <- mod_245.get(0);
        mod_245.put(1, t);
    endrule
    rule rule_313;
        ChannelMessage t;
        t <- mod_213.get(0);
        mod_243.put(0, t);
    endrule
    rule rule_314;
        ChannelMessage t;
        t <- mod_215.get(0);
        mod_216.put(0, t);
    endrule
    rule rule_315;
        ChannelMessage t;
        t <- mod_228.get(0);
        mod_227.put(0, t);
    endrule
    rule rule_316;
        ChannelMessage t;
        t <- mod_236.get(0);
        mod_235.put(0, t);
    endrule
    rule rule_317;
        ChannelMessage t;
        t <- mod_209.get(1);
        mod_210.put(0, t);
    endrule
    rule rule_318;
        ChannelMessage t;
        t <- mod_234.get(0);
        mod_233.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_206.put(0, t);
        end
        if (i == 1) begin
            mod_222.put(0, t);
        end
        if (i == 2) begin
            mod_228.put(0, t);
        end
        if (i == 3) begin
            mod_236.put(0, t);
        end
        if (i == 4) begin
            mod_242.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_210.get(0);
        end
        if (i == 2) begin
            t <- mod_210.get(1);
        end
        if (i == 0) begin
            t <- mod_210.get(2);
        end
        if (i == 3) begin
            t <- mod_222.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6040 (Operation_IFC);
    Operation_IFC mod_247_inner <- mkReshape(2, 64);
    Operation_IFC mod_247 <- mkDebugOperation(mod_247_inner, "mod_247");
    Operation_IFC mod_248_inner <- mkFlatten(1);
    Operation_IFC mod_248 <- mkDebugOperation(mod_248_inner, "mod_248");
    Operation_IFC mod_249_inner <- mkFlatten(2);
    Operation_IFC mod_249 <- mkDebugOperation(mod_249_inner, "mod_249");
    Operation_IFC mod_250_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_250 <- mkDebugOperation(mod_250_inner, "mod_250");
    Broadcast_IFC#(4) mod_251_inner <- mkBroadcast(4);
    Operation_IFC mod_251 <- mkDebugOperation(mod_251_inner.op, "mod_251");
    PMU_IFC mod_252_bufferize <- mkPMU(2);
    Operation_IFC mod_252_inner = mod_252_bufferize.operation;
    Operation_IFC mod_252 <- mkDebugOperation(mod_252_inner, "mod_252");
    Broadcast_IFC#(2) mod_253_inner <- mkBroadcast(2);
    Operation_IFC mod_253 <- mkDebugOperation(mod_253_inner.op, "mod_253");
    PMU_IFC mod_254_bufferize <- mkPMU(1);
    Operation_IFC mod_254_inner = mod_254_bufferize.operation;
    Operation_IFC mod_254 <- mkDebugOperation(mod_254_inner, "mod_254");
    Operation_IFC mod_255_inner <- mkBinaryMap(1150, matmul_t_tile);
    Operation_IFC mod_255 <- mkDebugOperation(mod_255_inner, "mod_255");
    Operation_IFC mod_256_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_256 <- mkDebugOperation(mod_256_inner, "mod_256");
    Operation_IFC mod_257_inner <- mkBinaryMap(1918, mul_tile);
    Operation_IFC mod_257 <- mkDebugOperation(mod_257_inner, "mod_257");
    PMU_IFC mod_258_bufferize <- mkPMU(1);
    Operation_IFC mod_258_inner = mod_258_bufferize.operation;
    Operation_IFC mod_258 <- mkDebugOperation(mod_258_inner, "mod_258");
    Operation_IFC mod_259_inner <- mkBinaryMap(2551, matmul_t_tile);
    Operation_IFC mod_259 <- mkDebugOperation(mod_259_inner, "mod_259");
    Operation_IFC mod_260_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_260 <- mkDebugOperation(mod_260_inner, "mod_260");
    Operation_IFC mod_261_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_261 <- mkDebugOperation(mod_261_inner, "mod_261");
    Operation_IFC mod_262_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_262 <- mkDebugOperation(mod_262_inner, "mod_262");
    Operation_IFC mod_263_inner <- mkBinaryMap(2817, mul_tile);
    Operation_IFC mod_263 <- mkDebugOperation(mod_263_inner, "mod_263");
    PMU_IFC mod_264_bufferize <- mkPMU(1);
    Operation_IFC mod_264_inner = mod_264_bufferize.operation;
    Operation_IFC mod_264 <- mkDebugOperation(mod_264_inner, "mod_264");
    PMU_IFC mod_265_bufferize <- mkPMU(2);
    Operation_IFC mod_265_inner = mod_265_bufferize.operation;
    Operation_IFC mod_265 <- mkDebugOperation(mod_265_inner, "mod_265");
    PMU_IFC mod_266_bufferize <- mkPMU(2);
    Operation_IFC mod_266_inner = mod_266_bufferize.operation;
    Operation_IFC mod_266 <- mkDebugOperation(mod_266_inner, "mod_266");
    Operation_IFC mod_267_inner <- mkRepeatStatic(8);
    Operation_IFC mod_267 <- mkDebugOperation(mod_267_inner, "mod_267");
    Operation_IFC mod_268_inner <- mkFlatten(1);
    Operation_IFC mod_268 <- mkDebugOperation(mod_268_inner, "mod_268");
    Operation_IFC mod_269_inner <- mkFlatten(0);
    Operation_IFC mod_269 <- mkDebugOperation(mod_269_inner, "mod_269");
    Operation_IFC mod_270_inner <- mkRepeatStatic(3);
    Operation_IFC mod_270 <- mkDebugOperation(mod_270_inner, "mod_270");
    Operation_IFC mod_271_inner <- mkUnaryMap(1790, silu_tile);
    Operation_IFC mod_271 <- mkDebugOperation(mod_271_inner, "mod_271");
    Operation_IFC mod_272_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_272 <- mkDebugOperation(mod_272_inner, "mod_272");
    Operation_IFC mod_273_inner <- mkBinaryMap(1662, matmul_t_tile);
    Operation_IFC mod_273 <- mkDebugOperation(mod_273_inner, "mod_273");
    PMU_IFC mod_274_bufferize <- mkPMU(2);
    Operation_IFC mod_274_inner = mod_274_bufferize.operation;
    Operation_IFC mod_274 <- mkDebugOperation(mod_274_inner, "mod_274");
    Operation_IFC mod_275_inner <- mkRepeatStatic(8);
    Operation_IFC mod_275 <- mkDebugOperation(mod_275_inner, "mod_275");
    Operation_IFC mod_276_inner <- mkFlatten(1);
    Operation_IFC mod_276 <- mkDebugOperation(mod_276_inner, "mod_276");
    Operation_IFC mod_277_inner <- mkFlatten(0);
    Operation_IFC mod_277 <- mkDebugOperation(mod_277_inner, "mod_277");
    PMU_IFC mod_278_bufferize <- mkPMU(1);
    Operation_IFC mod_278_inner = mod_278_bufferize.operation;
    Operation_IFC mod_278 <- mkDebugOperation(mod_278_inner, "mod_278");
    Operation_IFC mod_279_inner <- mkRepeatStatic(16);
    Operation_IFC mod_279 <- mkDebugOperation(mod_279_inner, "mod_279");
    PMU_IFC mod_280_bufferize <- mkPMU(2);
    Operation_IFC mod_280_inner = mod_280_bufferize.operation;
    Operation_IFC mod_280 <- mkDebugOperation(mod_280_inner, "mod_280");
    Operation_IFC mod_281_inner <- mkRepeatStatic(8);
    Operation_IFC mod_281 <- mkDebugOperation(mod_281_inner, "mod_281");
    Operation_IFC mod_282_inner <- mkFlatten(1);
    Operation_IFC mod_282 <- mkDebugOperation(mod_282_inner, "mod_282");
    Operation_IFC mod_283_inner <- mkFlatten(0);
    Operation_IFC mod_283 <- mkDebugOperation(mod_283_inner, "mod_283");
    Operation_IFC mod_284_inner <- mkRepeatStatic(16);
    Operation_IFC mod_284 <- mkDebugOperation(mod_284_inner, "mod_284");
    Operation_IFC mod_285_inner <- mkRepeatStatic(2);
    Operation_IFC mod_285 <- mkDebugOperation(mod_285_inner, "mod_285");
    PMU_IFC mod_286_bufferize <- mkPMU(2);
    Operation_IFC mod_286_inner = mod_286_bufferize.operation;
    Operation_IFC mod_286 <- mkDebugOperation(mod_286_inner, "mod_286");
    rule rule_319;
        ChannelMessage t;
        t <- mod_252.get(0);
        mod_285.put(0, t);
    endrule
    rule rule_320;
        ChannelMessage t;
        t <- mod_264.get(0);
        mod_264.put(1, t);
    endrule
    rule rule_321;
        ChannelMessage t;
        t <- mod_249.get(0);
        mod_250.put(0, t);
    endrule
    rule rule_322;
        ChannelMessage t;
        t <- mod_261.get(1);
        mod_262.put(0, t);
    endrule
    rule rule_323;
        ChannelMessage t;
        t <- mod_259.get(0);
        mod_260.put(0, t);
    endrule
    rule rule_324;
        ChannelMessage t;
        t <- mod_281.get(0);
        mod_280.put(1, t);
    endrule
    rule rule_325;
        ChannelMessage t;
        t <- mod_276.get(0);
        mod_274.put(0, t);
    endrule
    rule rule_326;
        ChannelMessage t;
        t <- mod_284.get(0);
        mod_254.put(1, t);
    endrule
    rule rule_327;
        ChannelMessage t;
        t <- mod_265.get(0);
        mod_265.put(1, t);
    endrule
    rule rule_328;
        ChannelMessage t;
        t <- mod_271.get(0);
        mod_257.put(1, t);
    endrule
    rule rule_329;
        ChannelMessage t;
        t <- mod_280.get(1);
        mod_255.put(1, t);
    endrule
    rule rule_330;
        ChannelMessage t;
        t <- mod_261.get(0);
        mod_265.put(0, t);
    endrule
    rule rule_331;
        ChannelMessage t;
        t <- mod_272.get(0);
        mod_271.put(0, t);
    endrule
    rule rule_332;
        ChannelMessage t;
        t <- mod_264.get(1);
        mod_262.put(1, t);
    endrule
    rule rule_333;
        ChannelMessage t;
        t <- mod_262.get(0);
        mod_264.put(0, t);
    endrule
    rule rule_334;
        ChannelMessage t;
        t <- mod_278.get(1);
        mod_273.put(0, t);
    endrule
    rule rule_335;
        ChannelMessage t;
        t <- mod_275.get(0);
        mod_274.put(1, t);
    endrule
    rule rule_336;
        ChannelMessage t;
        t <- mod_258.get(1);
        mod_259.put(0, t);
    endrule
    rule rule_337;
        ChannelMessage t;
        t <- mod_285.get(0);
        mod_252.put(1, t);
    endrule
    rule rule_338;
        ChannelMessage t;
        t <- mod_248.get(0);
        mod_249.put(0, t);
    endrule
    rule rule_339;
        ChannelMessage t;
        t <- mod_256.get(0);
        mod_257.put(0, t);
    endrule
    rule rule_340;
        ChannelMessage t;
        t <- mod_250.get(1);
        mod_251.put(0, t);
    endrule
    rule rule_341;
        ChannelMessage t;
        t <- mod_267.get(0);
        mod_266.put(1, t);
    endrule
    rule rule_342;
        ChannelMessage t;
        t <- mod_269.get(0);
        mod_268.put(0, t);
    endrule
    rule rule_343;
        ChannelMessage t;
        t <- mod_274.get(0);
        mod_275.put(0, t);
    endrule
    rule rule_344;
        ChannelMessage t;
        t <- mod_247.get(0);
        mod_248.put(0, t);
    endrule
    rule rule_345;
        ChannelMessage t;
        t <- mod_273.get(0);
        mod_272.put(0, t);
    endrule
    rule rule_346;
        ChannelMessage t;
        t <- mod_268.get(0);
        mod_266.put(0, t);
    endrule
    rule rule_347;
        ChannelMessage t;
        t <- mod_254.get(0);
        mod_284.put(0, t);
    endrule
    rule rule_348;
        ChannelMessage t;
        t <- mod_282.get(0);
        mod_280.put(0, t);
    endrule
    rule rule_349;
        ChannelMessage t;
        t <- mod_277.get(0);
        mod_276.put(0, t);
    endrule
    rule rule_350;
        ChannelMessage t;
        t <- mod_286.get(0);
        mod_286.put(1, t);
    endrule
    rule rule_351;
        ChannelMessage t;
        t <- mod_286.get(1);
        mod_250.put(1, t);
    endrule
    rule rule_352;
        ChannelMessage t;
        t <- mod_252.get(1);
        mod_253.put(0, t);
    endrule
    rule rule_353;
        ChannelMessage t;
        t <- mod_279.get(0);
        mod_278.put(1, t);
    endrule
    rule rule_354;
        ChannelMessage t;
        t <- mod_260.get(0);
        mod_261.put(0, t);
    endrule
    rule rule_355;
        ChannelMessage t;
        t <- mod_250.get(0);
        mod_286.put(0, t);
    endrule
    rule rule_356;
        ChannelMessage t;
        t <- mod_253.get(1);
        mod_254.put(0, t);
    endrule
    rule rule_357;
        ChannelMessage t;
        t <- mod_274.get(1);
        mod_273.put(1, t);
    endrule
    rule rule_358;
        ChannelMessage t;
        t <- mod_280.get(0);
        mod_281.put(0, t);
    endrule
    rule rule_359;
        ChannelMessage t;
        t <- mod_262.get(1);
        mod_263.put(1, t);
    endrule
    rule rule_360;
        ChannelMessage t;
        t <- mod_265.get(1);
        mod_261.put(1, t);
    endrule
    rule rule_361;
        ChannelMessage t;
        t <- mod_251.get(3);
        mod_252.put(0, t);
    endrule
    rule rule_362;
        ChannelMessage t;
        t <- mod_257.get(0);
        mod_258.put(0, t);
    endrule
    rule rule_363;
        ChannelMessage t;
        t <- mod_255.get(0);
        mod_256.put(0, t);
    endrule
    rule rule_364;
        ChannelMessage t;
        t <- mod_266.get(0);
        mod_267.put(0, t);
    endrule
    rule rule_365;
        ChannelMessage t;
        t <- mod_266.get(1);
        mod_259.put(1, t);
    endrule
    rule rule_366;
        ChannelMessage t;
        t <- mod_253.get(0);
        mod_278.put(0, t);
    endrule
    rule rule_367;
        ChannelMessage t;
        t <- mod_270.get(0);
        mod_258.put(1, t);
    endrule
    rule rule_368;
        ChannelMessage t;
        t <- mod_278.get(0);
        mod_279.put(0, t);
    endrule
    rule rule_369;
        ChannelMessage t;
        t <- mod_283.get(0);
        mod_282.put(0, t);
    endrule
    rule rule_370;
        ChannelMessage t;
        t <- mod_254.get(1);
        mod_255.put(0, t);
    endrule
    rule rule_371;
        ChannelMessage t;
        t <- mod_258.get(0);
        mod_270.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_247.put(0, t);
        end
        if (i == 1) begin
            mod_263.put(0, t);
        end
        if (i == 2) begin
            mod_269.put(0, t);
        end
        if (i == 3) begin
            mod_277.put(0, t);
        end
        if (i == 4) begin
            mod_283.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_251.get(0);
        end
        if (i == 1) begin
            t <- mod_251.get(1);
        end
        if (i == 3) begin
            t <- mod_251.get(2);
        end
        if (i == 2) begin
            t <- mod_263.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6041 (Operation_IFC);
    Operation_IFC mod_288_inner <- mkReshape(2, 64);
    Operation_IFC mod_288 <- mkDebugOperation(mod_288_inner, "mod_288");
    Operation_IFC mod_289_inner <- mkFlatten(1);
    Operation_IFC mod_289 <- mkDebugOperation(mod_289_inner, "mod_289");
    Operation_IFC mod_290_inner <- mkFlatten(2);
    Operation_IFC mod_290 <- mkDebugOperation(mod_290_inner, "mod_290");
    Operation_IFC mod_291_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_291 <- mkDebugOperation(mod_291_inner, "mod_291");
    Broadcast_IFC#(4) mod_292_inner <- mkBroadcast(4);
    Operation_IFC mod_292 <- mkDebugOperation(mod_292_inner.op, "mod_292");
    PMU_IFC mod_293_bufferize <- mkPMU(2);
    Operation_IFC mod_293_inner = mod_293_bufferize.operation;
    Operation_IFC mod_293 <- mkDebugOperation(mod_293_inner, "mod_293");
    Broadcast_IFC#(2) mod_294_inner <- mkBroadcast(2);
    Operation_IFC mod_294 <- mkDebugOperation(mod_294_inner.op, "mod_294");
    PMU_IFC mod_295_bufferize <- mkPMU(1);
    Operation_IFC mod_295_inner = mod_295_bufferize.operation;
    Operation_IFC mod_295 <- mkDebugOperation(mod_295_inner, "mod_295");
    Operation_IFC mod_296_inner <- mkBinaryMap(1149, matmul_t_tile);
    Operation_IFC mod_296 <- mkDebugOperation(mod_296_inner, "mod_296");
    Operation_IFC mod_297_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_297 <- mkDebugOperation(mod_297_inner, "mod_297");
    Operation_IFC mod_298_inner <- mkBinaryMap(1917, mul_tile);
    Operation_IFC mod_298 <- mkDebugOperation(mod_298_inner, "mod_298");
    PMU_IFC mod_299_bufferize <- mkPMU(1);
    Operation_IFC mod_299_inner = mod_299_bufferize.operation;
    Operation_IFC mod_299 <- mkDebugOperation(mod_299_inner, "mod_299");
    Operation_IFC mod_300_inner <- mkBinaryMap(2549, matmul_t_tile);
    Operation_IFC mod_300 <- mkDebugOperation(mod_300_inner, "mod_300");
    Operation_IFC mod_301_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_301 <- mkDebugOperation(mod_301_inner, "mod_301");
    Operation_IFC mod_302_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_302 <- mkDebugOperation(mod_302_inner, "mod_302");
    Operation_IFC mod_303_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_303 <- mkDebugOperation(mod_303_inner, "mod_303");
    Operation_IFC mod_304_inner <- mkBinaryMap(2816, mul_tile);
    Operation_IFC mod_304 <- mkDebugOperation(mod_304_inner, "mod_304");
    PMU_IFC mod_305_bufferize <- mkPMU(1);
    Operation_IFC mod_305_inner = mod_305_bufferize.operation;
    Operation_IFC mod_305 <- mkDebugOperation(mod_305_inner, "mod_305");
    PMU_IFC mod_306_bufferize <- mkPMU(2);
    Operation_IFC mod_306_inner = mod_306_bufferize.operation;
    Operation_IFC mod_306 <- mkDebugOperation(mod_306_inner, "mod_306");
    PMU_IFC mod_307_bufferize <- mkPMU(2);
    Operation_IFC mod_307_inner = mod_307_bufferize.operation;
    Operation_IFC mod_307 <- mkDebugOperation(mod_307_inner, "mod_307");
    Operation_IFC mod_308_inner <- mkRepeatStatic(8);
    Operation_IFC mod_308 <- mkDebugOperation(mod_308_inner, "mod_308");
    Operation_IFC mod_309_inner <- mkFlatten(1);
    Operation_IFC mod_309 <- mkDebugOperation(mod_309_inner, "mod_309");
    Operation_IFC mod_310_inner <- mkFlatten(0);
    Operation_IFC mod_310 <- mkDebugOperation(mod_310_inner, "mod_310");
    Operation_IFC mod_311_inner <- mkRepeatStatic(3);
    Operation_IFC mod_311 <- mkDebugOperation(mod_311_inner, "mod_311");
    Operation_IFC mod_312_inner <- mkUnaryMap(1789, silu_tile);
    Operation_IFC mod_312 <- mkDebugOperation(mod_312_inner, "mod_312");
    Operation_IFC mod_313_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_313 <- mkDebugOperation(mod_313_inner, "mod_313");
    Operation_IFC mod_314_inner <- mkBinaryMap(1661, matmul_t_tile);
    Operation_IFC mod_314 <- mkDebugOperation(mod_314_inner, "mod_314");
    PMU_IFC mod_315_bufferize <- mkPMU(2);
    Operation_IFC mod_315_inner = mod_315_bufferize.operation;
    Operation_IFC mod_315 <- mkDebugOperation(mod_315_inner, "mod_315");
    Operation_IFC mod_316_inner <- mkRepeatStatic(8);
    Operation_IFC mod_316 <- mkDebugOperation(mod_316_inner, "mod_316");
    Operation_IFC mod_317_inner <- mkFlatten(1);
    Operation_IFC mod_317 <- mkDebugOperation(mod_317_inner, "mod_317");
    Operation_IFC mod_318_inner <- mkFlatten(0);
    Operation_IFC mod_318 <- mkDebugOperation(mod_318_inner, "mod_318");
    PMU_IFC mod_319_bufferize <- mkPMU(1);
    Operation_IFC mod_319_inner = mod_319_bufferize.operation;
    Operation_IFC mod_319 <- mkDebugOperation(mod_319_inner, "mod_319");
    Operation_IFC mod_320_inner <- mkRepeatStatic(16);
    Operation_IFC mod_320 <- mkDebugOperation(mod_320_inner, "mod_320");
    PMU_IFC mod_321_bufferize <- mkPMU(2);
    Operation_IFC mod_321_inner = mod_321_bufferize.operation;
    Operation_IFC mod_321 <- mkDebugOperation(mod_321_inner, "mod_321");
    Operation_IFC mod_322_inner <- mkRepeatStatic(8);
    Operation_IFC mod_322 <- mkDebugOperation(mod_322_inner, "mod_322");
    Operation_IFC mod_323_inner <- mkFlatten(1);
    Operation_IFC mod_323 <- mkDebugOperation(mod_323_inner, "mod_323");
    Operation_IFC mod_324_inner <- mkFlatten(0);
    Operation_IFC mod_324 <- mkDebugOperation(mod_324_inner, "mod_324");
    Operation_IFC mod_325_inner <- mkRepeatStatic(16);
    Operation_IFC mod_325 <- mkDebugOperation(mod_325_inner, "mod_325");
    Operation_IFC mod_326_inner <- mkRepeatStatic(2);
    Operation_IFC mod_326 <- mkDebugOperation(mod_326_inner, "mod_326");
    PMU_IFC mod_327_bufferize <- mkPMU(2);
    Operation_IFC mod_327_inner = mod_327_bufferize.operation;
    Operation_IFC mod_327 <- mkDebugOperation(mod_327_inner, "mod_327");
    rule rule_372;
        ChannelMessage t;
        t <- mod_309.get(0);
        mod_307.put(0, t);
    endrule
    rule rule_373;
        ChannelMessage t;
        t <- mod_290.get(0);
        mod_291.put(0, t);
    endrule
    rule rule_374;
        ChannelMessage t;
        t <- mod_300.get(0);
        mod_301.put(0, t);
    endrule
    rule rule_375;
        ChannelMessage t;
        t <- mod_293.get(0);
        mod_326.put(0, t);
    endrule
    rule rule_376;
        ChannelMessage t;
        t <- mod_327.get(0);
        mod_327.put(1, t);
    endrule
    rule rule_377;
        ChannelMessage t;
        t <- mod_303.get(1);
        mod_304.put(1, t);
    endrule
    rule rule_378;
        ChannelMessage t;
        t <- mod_305.get(1);
        mod_303.put(1, t);
    endrule
    rule rule_379;
        ChannelMessage t;
        t <- mod_291.get(1);
        mod_292.put(0, t);
    endrule
    rule rule_380;
        ChannelMessage t;
        t <- mod_297.get(0);
        mod_298.put(0, t);
    endrule
    rule rule_381;
        ChannelMessage t;
        t <- mod_315.get(1);
        mod_314.put(1, t);
    endrule
    rule rule_382;
        ChannelMessage t;
        t <- mod_292.get(3);
        mod_293.put(0, t);
    endrule
    rule rule_383;
        ChannelMessage t;
        t <- mod_305.get(0);
        mod_305.put(1, t);
    endrule
    rule rule_384;
        ChannelMessage t;
        t <- mod_295.get(1);
        mod_296.put(0, t);
    endrule
    rule rule_385;
        ChannelMessage t;
        t <- mod_307.get(1);
        mod_300.put(1, t);
    endrule
    rule rule_386;
        ChannelMessage t;
        t <- mod_325.get(0);
        mod_295.put(1, t);
    endrule
    rule rule_387;
        ChannelMessage t;
        t <- mod_306.get(1);
        mod_302.put(1, t);
    endrule
    rule rule_388;
        ChannelMessage t;
        t <- mod_324.get(0);
        mod_323.put(0, t);
    endrule
    rule rule_389;
        ChannelMessage t;
        t <- mod_298.get(0);
        mod_299.put(0, t);
    endrule
    rule rule_390;
        ChannelMessage t;
        t <- mod_291.get(0);
        mod_327.put(0, t);
    endrule
    rule rule_391;
        ChannelMessage t;
        t <- mod_320.get(0);
        mod_319.put(1, t);
    endrule
    rule rule_392;
        ChannelMessage t;
        t <- mod_302.get(0);
        mod_306.put(0, t);
    endrule
    rule rule_393;
        ChannelMessage t;
        t <- mod_306.get(0);
        mod_306.put(1, t);
    endrule
    rule rule_394;
        ChannelMessage t;
        t <- mod_294.get(0);
        mod_319.put(0, t);
    endrule
    rule rule_395;
        ChannelMessage t;
        t <- mod_289.get(0);
        mod_290.put(0, t);
    endrule
    rule rule_396;
        ChannelMessage t;
        t <- mod_321.get(1);
        mod_296.put(1, t);
    endrule
    rule rule_397;
        ChannelMessage t;
        t <- mod_315.get(0);
        mod_316.put(0, t);
    endrule
    rule rule_398;
        ChannelMessage t;
        t <- mod_295.get(0);
        mod_325.put(0, t);
    endrule
    rule rule_399;
        ChannelMessage t;
        t <- mod_294.get(1);
        mod_295.put(0, t);
    endrule
    rule rule_400;
        ChannelMessage t;
        t <- mod_310.get(0);
        mod_309.put(0, t);
    endrule
    rule rule_401;
        ChannelMessage t;
        t <- mod_319.get(1);
        mod_314.put(0, t);
    endrule
    rule rule_402;
        ChannelMessage t;
        t <- mod_313.get(0);
        mod_312.put(0, t);
    endrule
    rule rule_403;
        ChannelMessage t;
        t <- mod_323.get(0);
        mod_321.put(0, t);
    endrule
    rule rule_404;
        ChannelMessage t;
        t <- mod_317.get(0);
        mod_315.put(0, t);
    endrule
    rule rule_405;
        ChannelMessage t;
        t <- mod_327.get(1);
        mod_291.put(1, t);
    endrule
    rule rule_406;
        ChannelMessage t;
        t <- mod_288.get(0);
        mod_289.put(0, t);
    endrule
    rule rule_407;
        ChannelMessage t;
        t <- mod_312.get(0);
        mod_298.put(1, t);
    endrule
    rule rule_408;
        ChannelMessage t;
        t <- mod_301.get(0);
        mod_302.put(0, t);
    endrule
    rule rule_409;
        ChannelMessage t;
        t <- mod_307.get(0);
        mod_308.put(0, t);
    endrule
    rule rule_410;
        ChannelMessage t;
        t <- mod_311.get(0);
        mod_299.put(1, t);
    endrule
    rule rule_411;
        ChannelMessage t;
        t <- mod_316.get(0);
        mod_315.put(1, t);
    endrule
    rule rule_412;
        ChannelMessage t;
        t <- mod_308.get(0);
        mod_307.put(1, t);
    endrule
    rule rule_413;
        ChannelMessage t;
        t <- mod_319.get(0);
        mod_320.put(0, t);
    endrule
    rule rule_414;
        ChannelMessage t;
        t <- mod_293.get(1);
        mod_294.put(0, t);
    endrule
    rule rule_415;
        ChannelMessage t;
        t <- mod_299.get(0);
        mod_311.put(0, t);
    endrule
    rule rule_416;
        ChannelMessage t;
        t <- mod_318.get(0);
        mod_317.put(0, t);
    endrule
    rule rule_417;
        ChannelMessage t;
        t <- mod_321.get(0);
        mod_322.put(0, t);
    endrule
    rule rule_418;
        ChannelMessage t;
        t <- mod_303.get(0);
        mod_305.put(0, t);
    endrule
    rule rule_419;
        ChannelMessage t;
        t <- mod_296.get(0);
        mod_297.put(0, t);
    endrule
    rule rule_420;
        ChannelMessage t;
        t <- mod_326.get(0);
        mod_293.put(1, t);
    endrule
    rule rule_421;
        ChannelMessage t;
        t <- mod_322.get(0);
        mod_321.put(1, t);
    endrule
    rule rule_422;
        ChannelMessage t;
        t <- mod_302.get(1);
        mod_303.put(0, t);
    endrule
    rule rule_423;
        ChannelMessage t;
        t <- mod_299.get(1);
        mod_300.put(0, t);
    endrule
    rule rule_424;
        ChannelMessage t;
        t <- mod_314.get(0);
        mod_313.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_288.put(0, t);
        end
        if (i == 1) begin
            mod_304.put(0, t);
        end
        if (i == 2) begin
            mod_310.put(0, t);
        end
        if (i == 3) begin
            mod_318.put(0, t);
        end
        if (i == 4) begin
            mod_324.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_292.get(0);
        end
        if (i == 3) begin
            t <- mod_292.get(1);
        end
        if (i == 1) begin
            t <- mod_292.get(2);
        end
        if (i == 2) begin
            t <- mod_304.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6042 (Operation_IFC);
    Operation_IFC mod_329_inner <- mkReshape(2, 64);
    Operation_IFC mod_329 <- mkDebugOperation(mod_329_inner, "mod_329");
    Operation_IFC mod_330_inner <- mkFlatten(1);
    Operation_IFC mod_330 <- mkDebugOperation(mod_330_inner, "mod_330");
    Operation_IFC mod_331_inner <- mkFlatten(2);
    Operation_IFC mod_331 <- mkDebugOperation(mod_331_inner, "mod_331");
    Operation_IFC mod_332_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_332 <- mkDebugOperation(mod_332_inner, "mod_332");
    Broadcast_IFC#(4) mod_333_inner <- mkBroadcast(4);
    Operation_IFC mod_333 <- mkDebugOperation(mod_333_inner.op, "mod_333");
    PMU_IFC mod_334_bufferize <- mkPMU(2);
    Operation_IFC mod_334_inner = mod_334_bufferize.operation;
    Operation_IFC mod_334 <- mkDebugOperation(mod_334_inner, "mod_334");
    Broadcast_IFC#(2) mod_335_inner <- mkBroadcast(2);
    Operation_IFC mod_335 <- mkDebugOperation(mod_335_inner.op, "mod_335");
    PMU_IFC mod_336_bufferize <- mkPMU(1);
    Operation_IFC mod_336_inner = mod_336_bufferize.operation;
    Operation_IFC mod_336 <- mkDebugOperation(mod_336_inner, "mod_336");
    Operation_IFC mod_337_inner <- mkBinaryMap(1148, matmul_t_tile);
    Operation_IFC mod_337 <- mkDebugOperation(mod_337_inner, "mod_337");
    Operation_IFC mod_338_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_338 <- mkDebugOperation(mod_338_inner, "mod_338");
    Operation_IFC mod_339_inner <- mkBinaryMap(1916, mul_tile);
    Operation_IFC mod_339 <- mkDebugOperation(mod_339_inner, "mod_339");
    PMU_IFC mod_340_bufferize <- mkPMU(1);
    Operation_IFC mod_340_inner = mod_340_bufferize.operation;
    Operation_IFC mod_340 <- mkDebugOperation(mod_340_inner, "mod_340");
    Operation_IFC mod_341_inner <- mkBinaryMap(2547, matmul_t_tile);
    Operation_IFC mod_341 <- mkDebugOperation(mod_341_inner, "mod_341");
    Operation_IFC mod_342_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_342 <- mkDebugOperation(mod_342_inner, "mod_342");
    Operation_IFC mod_343_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_343 <- mkDebugOperation(mod_343_inner, "mod_343");
    Operation_IFC mod_344_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_344 <- mkDebugOperation(mod_344_inner, "mod_344");
    Operation_IFC mod_345_inner <- mkBinaryMap(2815, mul_tile);
    Operation_IFC mod_345 <- mkDebugOperation(mod_345_inner, "mod_345");
    PMU_IFC mod_346_bufferize <- mkPMU(1);
    Operation_IFC mod_346_inner = mod_346_bufferize.operation;
    Operation_IFC mod_346 <- mkDebugOperation(mod_346_inner, "mod_346");
    PMU_IFC mod_347_bufferize <- mkPMU(2);
    Operation_IFC mod_347_inner = mod_347_bufferize.operation;
    Operation_IFC mod_347 <- mkDebugOperation(mod_347_inner, "mod_347");
    PMU_IFC mod_348_bufferize <- mkPMU(2);
    Operation_IFC mod_348_inner = mod_348_bufferize.operation;
    Operation_IFC mod_348 <- mkDebugOperation(mod_348_inner, "mod_348");
    Operation_IFC mod_349_inner <- mkRepeatStatic(8);
    Operation_IFC mod_349 <- mkDebugOperation(mod_349_inner, "mod_349");
    Operation_IFC mod_350_inner <- mkFlatten(1);
    Operation_IFC mod_350 <- mkDebugOperation(mod_350_inner, "mod_350");
    Operation_IFC mod_351_inner <- mkFlatten(0);
    Operation_IFC mod_351 <- mkDebugOperation(mod_351_inner, "mod_351");
    Operation_IFC mod_352_inner <- mkRepeatStatic(3);
    Operation_IFC mod_352 <- mkDebugOperation(mod_352_inner, "mod_352");
    Operation_IFC mod_353_inner <- mkUnaryMap(1788, silu_tile);
    Operation_IFC mod_353 <- mkDebugOperation(mod_353_inner, "mod_353");
    Operation_IFC mod_354_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_354 <- mkDebugOperation(mod_354_inner, "mod_354");
    Operation_IFC mod_355_inner <- mkBinaryMap(1660, matmul_t_tile);
    Operation_IFC mod_355 <- mkDebugOperation(mod_355_inner, "mod_355");
    PMU_IFC mod_356_bufferize <- mkPMU(2);
    Operation_IFC mod_356_inner = mod_356_bufferize.operation;
    Operation_IFC mod_356 <- mkDebugOperation(mod_356_inner, "mod_356");
    Operation_IFC mod_357_inner <- mkRepeatStatic(8);
    Operation_IFC mod_357 <- mkDebugOperation(mod_357_inner, "mod_357");
    Operation_IFC mod_358_inner <- mkFlatten(1);
    Operation_IFC mod_358 <- mkDebugOperation(mod_358_inner, "mod_358");
    Operation_IFC mod_359_inner <- mkFlatten(0);
    Operation_IFC mod_359 <- mkDebugOperation(mod_359_inner, "mod_359");
    PMU_IFC mod_360_bufferize <- mkPMU(1);
    Operation_IFC mod_360_inner = mod_360_bufferize.operation;
    Operation_IFC mod_360 <- mkDebugOperation(mod_360_inner, "mod_360");
    Operation_IFC mod_361_inner <- mkRepeatStatic(16);
    Operation_IFC mod_361 <- mkDebugOperation(mod_361_inner, "mod_361");
    PMU_IFC mod_362_bufferize <- mkPMU(2);
    Operation_IFC mod_362_inner = mod_362_bufferize.operation;
    Operation_IFC mod_362 <- mkDebugOperation(mod_362_inner, "mod_362");
    Operation_IFC mod_363_inner <- mkRepeatStatic(8);
    Operation_IFC mod_363 <- mkDebugOperation(mod_363_inner, "mod_363");
    Operation_IFC mod_364_inner <- mkFlatten(1);
    Operation_IFC mod_364 <- mkDebugOperation(mod_364_inner, "mod_364");
    Operation_IFC mod_365_inner <- mkFlatten(0);
    Operation_IFC mod_365 <- mkDebugOperation(mod_365_inner, "mod_365");
    Operation_IFC mod_366_inner <- mkRepeatStatic(16);
    Operation_IFC mod_366 <- mkDebugOperation(mod_366_inner, "mod_366");
    Operation_IFC mod_367_inner <- mkRepeatStatic(2);
    Operation_IFC mod_367 <- mkDebugOperation(mod_367_inner, "mod_367");
    PMU_IFC mod_368_bufferize <- mkPMU(2);
    Operation_IFC mod_368_inner = mod_368_bufferize.operation;
    Operation_IFC mod_368 <- mkDebugOperation(mod_368_inner, "mod_368");
    rule rule_425;
        ChannelMessage t;
        t <- mod_368.get(1);
        mod_332.put(1, t);
    endrule
    rule rule_426;
        ChannelMessage t;
        t <- mod_334.get(1);
        mod_335.put(0, t);
    endrule
    rule rule_427;
        ChannelMessage t;
        t <- mod_351.get(0);
        mod_350.put(0, t);
    endrule
    rule rule_428;
        ChannelMessage t;
        t <- mod_342.get(0);
        mod_343.put(0, t);
    endrule
    rule rule_429;
        ChannelMessage t;
        t <- mod_360.get(1);
        mod_355.put(0, t);
    endrule
    rule rule_430;
        ChannelMessage t;
        t <- mod_338.get(0);
        mod_339.put(0, t);
    endrule
    rule rule_431;
        ChannelMessage t;
        t <- mod_330.get(0);
        mod_331.put(0, t);
    endrule
    rule rule_432;
        ChannelMessage t;
        t <- mod_365.get(0);
        mod_364.put(0, t);
    endrule
    rule rule_433;
        ChannelMessage t;
        t <- mod_346.get(0);
        mod_346.put(1, t);
    endrule
    rule rule_434;
        ChannelMessage t;
        t <- mod_353.get(0);
        mod_339.put(1, t);
    endrule
    rule rule_435;
        ChannelMessage t;
        t <- mod_359.get(0);
        mod_358.put(0, t);
    endrule
    rule rule_436;
        ChannelMessage t;
        t <- mod_360.get(0);
        mod_361.put(0, t);
    endrule
    rule rule_437;
        ChannelMessage t;
        t <- mod_352.get(0);
        mod_340.put(1, t);
    endrule
    rule rule_438;
        ChannelMessage t;
        t <- mod_356.get(1);
        mod_355.put(1, t);
    endrule
    rule rule_439;
        ChannelMessage t;
        t <- mod_341.get(0);
        mod_342.put(0, t);
    endrule
    rule rule_440;
        ChannelMessage t;
        t <- mod_340.get(1);
        mod_341.put(0, t);
    endrule
    rule rule_441;
        ChannelMessage t;
        t <- mod_367.get(0);
        mod_334.put(1, t);
    endrule
    rule rule_442;
        ChannelMessage t;
        t <- mod_358.get(0);
        mod_356.put(0, t);
    endrule
    rule rule_443;
        ChannelMessage t;
        t <- mod_333.get(3);
        mod_334.put(0, t);
    endrule
    rule rule_444;
        ChannelMessage t;
        t <- mod_348.get(1);
        mod_341.put(1, t);
    endrule
    rule rule_445;
        ChannelMessage t;
        t <- mod_357.get(0);
        mod_356.put(1, t);
    endrule
    rule rule_446;
        ChannelMessage t;
        t <- mod_335.get(1);
        mod_336.put(0, t);
    endrule
    rule rule_447;
        ChannelMessage t;
        t <- mod_336.get(1);
        mod_337.put(0, t);
    endrule
    rule rule_448;
        ChannelMessage t;
        t <- mod_340.get(0);
        mod_352.put(0, t);
    endrule
    rule rule_449;
        ChannelMessage t;
        t <- mod_335.get(0);
        mod_360.put(0, t);
    endrule
    rule rule_450;
        ChannelMessage t;
        t <- mod_349.get(0);
        mod_348.put(1, t);
    endrule
    rule rule_451;
        ChannelMessage t;
        t <- mod_332.get(0);
        mod_368.put(0, t);
    endrule
    rule rule_452;
        ChannelMessage t;
        t <- mod_337.get(0);
        mod_338.put(0, t);
    endrule
    rule rule_453;
        ChannelMessage t;
        t <- mod_343.get(0);
        mod_347.put(0, t);
    endrule
    rule rule_454;
        ChannelMessage t;
        t <- mod_356.get(0);
        mod_357.put(0, t);
    endrule
    rule rule_455;
        ChannelMessage t;
        t <- mod_366.get(0);
        mod_336.put(1, t);
    endrule
    rule rule_456;
        ChannelMessage t;
        t <- mod_346.get(1);
        mod_344.put(1, t);
    endrule
    rule rule_457;
        ChannelMessage t;
        t <- mod_362.get(0);
        mod_363.put(0, t);
    endrule
    rule rule_458;
        ChannelMessage t;
        t <- mod_336.get(0);
        mod_366.put(0, t);
    endrule
    rule rule_459;
        ChannelMessage t;
        t <- mod_350.get(0);
        mod_348.put(0, t);
    endrule
    rule rule_460;
        ChannelMessage t;
        t <- mod_331.get(0);
        mod_332.put(0, t);
    endrule
    rule rule_461;
        ChannelMessage t;
        t <- mod_364.get(0);
        mod_362.put(0, t);
    endrule
    rule rule_462;
        ChannelMessage t;
        t <- mod_354.get(0);
        mod_353.put(0, t);
    endrule
    rule rule_463;
        ChannelMessage t;
        t <- mod_329.get(0);
        mod_330.put(0, t);
    endrule
    rule rule_464;
        ChannelMessage t;
        t <- mod_339.get(0);
        mod_340.put(0, t);
    endrule
    rule rule_465;
        ChannelMessage t;
        t <- mod_361.get(0);
        mod_360.put(1, t);
    endrule
    rule rule_466;
        ChannelMessage t;
        t <- mod_347.get(0);
        mod_347.put(1, t);
    endrule
    rule rule_467;
        ChannelMessage t;
        t <- mod_347.get(1);
        mod_343.put(1, t);
    endrule
    rule rule_468;
        ChannelMessage t;
        t <- mod_332.get(1);
        mod_333.put(0, t);
    endrule
    rule rule_469;
        ChannelMessage t;
        t <- mod_363.get(0);
        mod_362.put(1, t);
    endrule
    rule rule_470;
        ChannelMessage t;
        t <- mod_348.get(0);
        mod_349.put(0, t);
    endrule
    rule rule_471;
        ChannelMessage t;
        t <- mod_355.get(0);
        mod_354.put(0, t);
    endrule
    rule rule_472;
        ChannelMessage t;
        t <- mod_344.get(0);
        mod_346.put(0, t);
    endrule
    rule rule_473;
        ChannelMessage t;
        t <- mod_368.get(0);
        mod_368.put(1, t);
    endrule
    rule rule_474;
        ChannelMessage t;
        t <- mod_344.get(1);
        mod_345.put(1, t);
    endrule
    rule rule_475;
        ChannelMessage t;
        t <- mod_334.get(0);
        mod_367.put(0, t);
    endrule
    rule rule_476;
        ChannelMessage t;
        t <- mod_343.get(1);
        mod_344.put(0, t);
    endrule
    rule rule_477;
        ChannelMessage t;
        t <- mod_362.get(1);
        mod_337.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_329.put(0, t);
        end
        if (i == 1) begin
            mod_345.put(0, t);
        end
        if (i == 2) begin
            mod_351.put(0, t);
        end
        if (i == 3) begin
            mod_359.put(0, t);
        end
        if (i == 4) begin
            mod_365.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_333.get(0);
        end
        if (i == 2) begin
            t <- mod_333.get(1);
        end
        if (i == 1) begin
            t <- mod_333.get(2);
        end
        if (i == 3) begin
            t <- mod_345.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6043 (Operation_IFC);
    Operation_IFC mod_370_inner <- mkReshape(2, 64);
    Operation_IFC mod_370 <- mkDebugOperation(mod_370_inner, "mod_370");
    Operation_IFC mod_371_inner <- mkFlatten(1);
    Operation_IFC mod_371 <- mkDebugOperation(mod_371_inner, "mod_371");
    Operation_IFC mod_372_inner <- mkFlatten(2);
    Operation_IFC mod_372 <- mkDebugOperation(mod_372_inner, "mod_372");
    Operation_IFC mod_373_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_373 <- mkDebugOperation(mod_373_inner, "mod_373");
    Broadcast_IFC#(4) mod_374_inner <- mkBroadcast(4);
    Operation_IFC mod_374 <- mkDebugOperation(mod_374_inner.op, "mod_374");
    PMU_IFC mod_375_bufferize <- mkPMU(2);
    Operation_IFC mod_375_inner = mod_375_bufferize.operation;
    Operation_IFC mod_375 <- mkDebugOperation(mod_375_inner, "mod_375");
    Broadcast_IFC#(2) mod_376_inner <- mkBroadcast(2);
    Operation_IFC mod_376 <- mkDebugOperation(mod_376_inner.op, "mod_376");
    PMU_IFC mod_377_bufferize <- mkPMU(1);
    Operation_IFC mod_377_inner = mod_377_bufferize.operation;
    Operation_IFC mod_377 <- mkDebugOperation(mod_377_inner, "mod_377");
    Operation_IFC mod_378_inner <- mkBinaryMap(1147, matmul_t_tile);
    Operation_IFC mod_378 <- mkDebugOperation(mod_378_inner, "mod_378");
    Operation_IFC mod_379_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_379 <- mkDebugOperation(mod_379_inner, "mod_379");
    Operation_IFC mod_380_inner <- mkBinaryMap(1915, mul_tile);
    Operation_IFC mod_380 <- mkDebugOperation(mod_380_inner, "mod_380");
    PMU_IFC mod_381_bufferize <- mkPMU(1);
    Operation_IFC mod_381_inner = mod_381_bufferize.operation;
    Operation_IFC mod_381 <- mkDebugOperation(mod_381_inner, "mod_381");
    Operation_IFC mod_382_inner <- mkBinaryMap(2545, matmul_t_tile);
    Operation_IFC mod_382 <- mkDebugOperation(mod_382_inner, "mod_382");
    Operation_IFC mod_383_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_383 <- mkDebugOperation(mod_383_inner, "mod_383");
    Operation_IFC mod_384_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_384 <- mkDebugOperation(mod_384_inner, "mod_384");
    Operation_IFC mod_385_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_385 <- mkDebugOperation(mod_385_inner, "mod_385");
    Operation_IFC mod_386_inner <- mkBinaryMap(2814, mul_tile);
    Operation_IFC mod_386 <- mkDebugOperation(mod_386_inner, "mod_386");
    PMU_IFC mod_387_bufferize <- mkPMU(1);
    Operation_IFC mod_387_inner = mod_387_bufferize.operation;
    Operation_IFC mod_387 <- mkDebugOperation(mod_387_inner, "mod_387");
    PMU_IFC mod_388_bufferize <- mkPMU(2);
    Operation_IFC mod_388_inner = mod_388_bufferize.operation;
    Operation_IFC mod_388 <- mkDebugOperation(mod_388_inner, "mod_388");
    PMU_IFC mod_389_bufferize <- mkPMU(2);
    Operation_IFC mod_389_inner = mod_389_bufferize.operation;
    Operation_IFC mod_389 <- mkDebugOperation(mod_389_inner, "mod_389");
    Operation_IFC mod_390_inner <- mkRepeatStatic(8);
    Operation_IFC mod_390 <- mkDebugOperation(mod_390_inner, "mod_390");
    Operation_IFC mod_391_inner <- mkFlatten(1);
    Operation_IFC mod_391 <- mkDebugOperation(mod_391_inner, "mod_391");
    Operation_IFC mod_392_inner <- mkFlatten(0);
    Operation_IFC mod_392 <- mkDebugOperation(mod_392_inner, "mod_392");
    Operation_IFC mod_393_inner <- mkRepeatStatic(3);
    Operation_IFC mod_393 <- mkDebugOperation(mod_393_inner, "mod_393");
    Operation_IFC mod_394_inner <- mkUnaryMap(1787, silu_tile);
    Operation_IFC mod_394 <- mkDebugOperation(mod_394_inner, "mod_394");
    Operation_IFC mod_395_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_395 <- mkDebugOperation(mod_395_inner, "mod_395");
    Operation_IFC mod_396_inner <- mkBinaryMap(1659, matmul_t_tile);
    Operation_IFC mod_396 <- mkDebugOperation(mod_396_inner, "mod_396");
    PMU_IFC mod_397_bufferize <- mkPMU(2);
    Operation_IFC mod_397_inner = mod_397_bufferize.operation;
    Operation_IFC mod_397 <- mkDebugOperation(mod_397_inner, "mod_397");
    Operation_IFC mod_398_inner <- mkRepeatStatic(8);
    Operation_IFC mod_398 <- mkDebugOperation(mod_398_inner, "mod_398");
    Operation_IFC mod_399_inner <- mkFlatten(1);
    Operation_IFC mod_399 <- mkDebugOperation(mod_399_inner, "mod_399");
    Operation_IFC mod_400_inner <- mkFlatten(0);
    Operation_IFC mod_400 <- mkDebugOperation(mod_400_inner, "mod_400");
    PMU_IFC mod_401_bufferize <- mkPMU(1);
    Operation_IFC mod_401_inner = mod_401_bufferize.operation;
    Operation_IFC mod_401 <- mkDebugOperation(mod_401_inner, "mod_401");
    Operation_IFC mod_402_inner <- mkRepeatStatic(16);
    Operation_IFC mod_402 <- mkDebugOperation(mod_402_inner, "mod_402");
    PMU_IFC mod_403_bufferize <- mkPMU(2);
    Operation_IFC mod_403_inner = mod_403_bufferize.operation;
    Operation_IFC mod_403 <- mkDebugOperation(mod_403_inner, "mod_403");
    Operation_IFC mod_404_inner <- mkRepeatStatic(8);
    Operation_IFC mod_404 <- mkDebugOperation(mod_404_inner, "mod_404");
    Operation_IFC mod_405_inner <- mkFlatten(1);
    Operation_IFC mod_405 <- mkDebugOperation(mod_405_inner, "mod_405");
    Operation_IFC mod_406_inner <- mkFlatten(0);
    Operation_IFC mod_406 <- mkDebugOperation(mod_406_inner, "mod_406");
    Operation_IFC mod_407_inner <- mkRepeatStatic(16);
    Operation_IFC mod_407 <- mkDebugOperation(mod_407_inner, "mod_407");
    Operation_IFC mod_408_inner <- mkRepeatStatic(2);
    Operation_IFC mod_408 <- mkDebugOperation(mod_408_inner, "mod_408");
    PMU_IFC mod_409_bufferize <- mkPMU(2);
    Operation_IFC mod_409_inner = mod_409_bufferize.operation;
    Operation_IFC mod_409 <- mkDebugOperation(mod_409_inner, "mod_409");
    rule rule_478;
        ChannelMessage t;
        t <- mod_382.get(0);
        mod_383.put(0, t);
    endrule
    rule rule_479;
        ChannelMessage t;
        t <- mod_401.get(0);
        mod_402.put(0, t);
    endrule
    rule rule_480;
        ChannelMessage t;
        t <- mod_407.get(0);
        mod_377.put(1, t);
    endrule
    rule rule_481;
        ChannelMessage t;
        t <- mod_383.get(0);
        mod_384.put(0, t);
    endrule
    rule rule_482;
        ChannelMessage t;
        t <- mod_375.get(0);
        mod_408.put(0, t);
    endrule
    rule rule_483;
        ChannelMessage t;
        t <- mod_397.get(1);
        mod_396.put(1, t);
    endrule
    rule rule_484;
        ChannelMessage t;
        t <- mod_405.get(0);
        mod_403.put(0, t);
    endrule
    rule rule_485;
        ChannelMessage t;
        t <- mod_389.get(1);
        mod_382.put(1, t);
    endrule
    rule rule_486;
        ChannelMessage t;
        t <- mod_376.get(0);
        mod_401.put(0, t);
    endrule
    rule rule_487;
        ChannelMessage t;
        t <- mod_397.get(0);
        mod_398.put(0, t);
    endrule
    rule rule_488;
        ChannelMessage t;
        t <- mod_377.get(0);
        mod_407.put(0, t);
    endrule
    rule rule_489;
        ChannelMessage t;
        t <- mod_402.get(0);
        mod_401.put(1, t);
    endrule
    rule rule_490;
        ChannelMessage t;
        t <- mod_385.get(0);
        mod_387.put(0, t);
    endrule
    rule rule_491;
        ChannelMessage t;
        t <- mod_403.get(0);
        mod_404.put(0, t);
    endrule
    rule rule_492;
        ChannelMessage t;
        t <- mod_390.get(0);
        mod_389.put(1, t);
    endrule
    rule rule_493;
        ChannelMessage t;
        t <- mod_378.get(0);
        mod_379.put(0, t);
    endrule
    rule rule_494;
        ChannelMessage t;
        t <- mod_381.get(1);
        mod_382.put(0, t);
    endrule
    rule rule_495;
        ChannelMessage t;
        t <- mod_387.get(1);
        mod_385.put(1, t);
    endrule
    rule rule_496;
        ChannelMessage t;
        t <- mod_399.get(0);
        mod_397.put(0, t);
    endrule
    rule rule_497;
        ChannelMessage t;
        t <- mod_373.get(0);
        mod_409.put(0, t);
    endrule
    rule rule_498;
        ChannelMessage t;
        t <- mod_392.get(0);
        mod_391.put(0, t);
    endrule
    rule rule_499;
        ChannelMessage t;
        t <- mod_404.get(0);
        mod_403.put(1, t);
    endrule
    rule rule_500;
        ChannelMessage t;
        t <- mod_388.get(0);
        mod_388.put(1, t);
    endrule
    rule rule_501;
        ChannelMessage t;
        t <- mod_375.get(1);
        mod_376.put(0, t);
    endrule
    rule rule_502;
        ChannelMessage t;
        t <- mod_409.get(0);
        mod_409.put(1, t);
    endrule
    rule rule_503;
        ChannelMessage t;
        t <- mod_373.get(1);
        mod_374.put(0, t);
    endrule
    rule rule_504;
        ChannelMessage t;
        t <- mod_376.get(1);
        mod_377.put(0, t);
    endrule
    rule rule_505;
        ChannelMessage t;
        t <- mod_381.get(0);
        mod_393.put(0, t);
    endrule
    rule rule_506;
        ChannelMessage t;
        t <- mod_377.get(1);
        mod_378.put(0, t);
    endrule
    rule rule_507;
        ChannelMessage t;
        t <- mod_391.get(0);
        mod_389.put(0, t);
    endrule
    rule rule_508;
        ChannelMessage t;
        t <- mod_394.get(0);
        mod_380.put(1, t);
    endrule
    rule rule_509;
        ChannelMessage t;
        t <- mod_389.get(0);
        mod_390.put(0, t);
    endrule
    rule rule_510;
        ChannelMessage t;
        t <- mod_396.get(0);
        mod_395.put(0, t);
    endrule
    rule rule_511;
        ChannelMessage t;
        t <- mod_403.get(1);
        mod_378.put(1, t);
    endrule
    rule rule_512;
        ChannelMessage t;
        t <- mod_401.get(1);
        mod_396.put(0, t);
    endrule
    rule rule_513;
        ChannelMessage t;
        t <- mod_406.get(0);
        mod_405.put(0, t);
    endrule
    rule rule_514;
        ChannelMessage t;
        t <- mod_384.get(1);
        mod_385.put(0, t);
    endrule
    rule rule_515;
        ChannelMessage t;
        t <- mod_409.get(1);
        mod_373.put(1, t);
    endrule
    rule rule_516;
        ChannelMessage t;
        t <- mod_370.get(0);
        mod_371.put(0, t);
    endrule
    rule rule_517;
        ChannelMessage t;
        t <- mod_371.get(0);
        mod_372.put(0, t);
    endrule
    rule rule_518;
        ChannelMessage t;
        t <- mod_374.get(3);
        mod_375.put(0, t);
    endrule
    rule rule_519;
        ChannelMessage t;
        t <- mod_379.get(0);
        mod_380.put(0, t);
    endrule
    rule rule_520;
        ChannelMessage t;
        t <- mod_408.get(0);
        mod_375.put(1, t);
    endrule
    rule rule_521;
        ChannelMessage t;
        t <- mod_380.get(0);
        mod_381.put(0, t);
    endrule
    rule rule_522;
        ChannelMessage t;
        t <- mod_372.get(0);
        mod_373.put(0, t);
    endrule
    rule rule_523;
        ChannelMessage t;
        t <- mod_395.get(0);
        mod_394.put(0, t);
    endrule
    rule rule_524;
        ChannelMessage t;
        t <- mod_388.get(1);
        mod_384.put(1, t);
    endrule
    rule rule_525;
        ChannelMessage t;
        t <- mod_384.get(0);
        mod_388.put(0, t);
    endrule
    rule rule_526;
        ChannelMessage t;
        t <- mod_387.get(0);
        mod_387.put(1, t);
    endrule
    rule rule_527;
        ChannelMessage t;
        t <- mod_398.get(0);
        mod_397.put(1, t);
    endrule
    rule rule_528;
        ChannelMessage t;
        t <- mod_385.get(1);
        mod_386.put(1, t);
    endrule
    rule rule_529;
        ChannelMessage t;
        t <- mod_393.get(0);
        mod_381.put(1, t);
    endrule
    rule rule_530;
        ChannelMessage t;
        t <- mod_400.get(0);
        mod_399.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_370.put(0, t);
        end
        if (i == 1) begin
            mod_386.put(0, t);
        end
        if (i == 2) begin
            mod_392.put(0, t);
        end
        if (i == 3) begin
            mod_400.put(0, t);
        end
        if (i == 4) begin
            mod_406.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_374.get(0);
        end
        if (i == 2) begin
            t <- mod_374.get(1);
        end
        if (i == 3) begin
            t <- mod_374.get(2);
        end
        if (i == 0) begin
            t <- mod_386.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6044 (Operation_IFC);
    Operation_IFC mod_411_inner <- mkReshape(2, 64);
    Operation_IFC mod_411 <- mkDebugOperation(mod_411_inner, "mod_411");
    Operation_IFC mod_412_inner <- mkFlatten(1);
    Operation_IFC mod_412 <- mkDebugOperation(mod_412_inner, "mod_412");
    Operation_IFC mod_413_inner <- mkFlatten(2);
    Operation_IFC mod_413 <- mkDebugOperation(mod_413_inner, "mod_413");
    Operation_IFC mod_414_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_414 <- mkDebugOperation(mod_414_inner, "mod_414");
    Broadcast_IFC#(4) mod_415_inner <- mkBroadcast(4);
    Operation_IFC mod_415 <- mkDebugOperation(mod_415_inner.op, "mod_415");
    PMU_IFC mod_416_bufferize <- mkPMU(2);
    Operation_IFC mod_416_inner = mod_416_bufferize.operation;
    Operation_IFC mod_416 <- mkDebugOperation(mod_416_inner, "mod_416");
    Broadcast_IFC#(2) mod_417_inner <- mkBroadcast(2);
    Operation_IFC mod_417 <- mkDebugOperation(mod_417_inner.op, "mod_417");
    PMU_IFC mod_418_bufferize <- mkPMU(1);
    Operation_IFC mod_418_inner = mod_418_bufferize.operation;
    Operation_IFC mod_418 <- mkDebugOperation(mod_418_inner, "mod_418");
    Operation_IFC mod_419_inner <- mkBinaryMap(1146, matmul_t_tile);
    Operation_IFC mod_419 <- mkDebugOperation(mod_419_inner, "mod_419");
    Operation_IFC mod_420_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_420 <- mkDebugOperation(mod_420_inner, "mod_420");
    Operation_IFC mod_421_inner <- mkBinaryMap(1914, mul_tile);
    Operation_IFC mod_421 <- mkDebugOperation(mod_421_inner, "mod_421");
    PMU_IFC mod_422_bufferize <- mkPMU(1);
    Operation_IFC mod_422_inner = mod_422_bufferize.operation;
    Operation_IFC mod_422 <- mkDebugOperation(mod_422_inner, "mod_422");
    Operation_IFC mod_423_inner <- mkBinaryMap(2543, matmul_t_tile);
    Operation_IFC mod_423 <- mkDebugOperation(mod_423_inner, "mod_423");
    Operation_IFC mod_424_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_424 <- mkDebugOperation(mod_424_inner, "mod_424");
    Operation_IFC mod_425_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_425 <- mkDebugOperation(mod_425_inner, "mod_425");
    Operation_IFC mod_426_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_426 <- mkDebugOperation(mod_426_inner, "mod_426");
    Operation_IFC mod_427_inner <- mkBinaryMap(2813, mul_tile);
    Operation_IFC mod_427 <- mkDebugOperation(mod_427_inner, "mod_427");
    PMU_IFC mod_428_bufferize <- mkPMU(1);
    Operation_IFC mod_428_inner = mod_428_bufferize.operation;
    Operation_IFC mod_428 <- mkDebugOperation(mod_428_inner, "mod_428");
    PMU_IFC mod_429_bufferize <- mkPMU(2);
    Operation_IFC mod_429_inner = mod_429_bufferize.operation;
    Operation_IFC mod_429 <- mkDebugOperation(mod_429_inner, "mod_429");
    PMU_IFC mod_430_bufferize <- mkPMU(2);
    Operation_IFC mod_430_inner = mod_430_bufferize.operation;
    Operation_IFC mod_430 <- mkDebugOperation(mod_430_inner, "mod_430");
    Operation_IFC mod_431_inner <- mkRepeatStatic(8);
    Operation_IFC mod_431 <- mkDebugOperation(mod_431_inner, "mod_431");
    Operation_IFC mod_432_inner <- mkFlatten(1);
    Operation_IFC mod_432 <- mkDebugOperation(mod_432_inner, "mod_432");
    Operation_IFC mod_433_inner <- mkFlatten(0);
    Operation_IFC mod_433 <- mkDebugOperation(mod_433_inner, "mod_433");
    Operation_IFC mod_434_inner <- mkRepeatStatic(3);
    Operation_IFC mod_434 <- mkDebugOperation(mod_434_inner, "mod_434");
    Operation_IFC mod_435_inner <- mkUnaryMap(1786, silu_tile);
    Operation_IFC mod_435 <- mkDebugOperation(mod_435_inner, "mod_435");
    Operation_IFC mod_436_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_436 <- mkDebugOperation(mod_436_inner, "mod_436");
    Operation_IFC mod_437_inner <- mkBinaryMap(1658, matmul_t_tile);
    Operation_IFC mod_437 <- mkDebugOperation(mod_437_inner, "mod_437");
    PMU_IFC mod_438_bufferize <- mkPMU(2);
    Operation_IFC mod_438_inner = mod_438_bufferize.operation;
    Operation_IFC mod_438 <- mkDebugOperation(mod_438_inner, "mod_438");
    Operation_IFC mod_439_inner <- mkRepeatStatic(8);
    Operation_IFC mod_439 <- mkDebugOperation(mod_439_inner, "mod_439");
    Operation_IFC mod_440_inner <- mkFlatten(1);
    Operation_IFC mod_440 <- mkDebugOperation(mod_440_inner, "mod_440");
    Operation_IFC mod_441_inner <- mkFlatten(0);
    Operation_IFC mod_441 <- mkDebugOperation(mod_441_inner, "mod_441");
    PMU_IFC mod_442_bufferize <- mkPMU(1);
    Operation_IFC mod_442_inner = mod_442_bufferize.operation;
    Operation_IFC mod_442 <- mkDebugOperation(mod_442_inner, "mod_442");
    Operation_IFC mod_443_inner <- mkRepeatStatic(16);
    Operation_IFC mod_443 <- mkDebugOperation(mod_443_inner, "mod_443");
    PMU_IFC mod_444_bufferize <- mkPMU(2);
    Operation_IFC mod_444_inner = mod_444_bufferize.operation;
    Operation_IFC mod_444 <- mkDebugOperation(mod_444_inner, "mod_444");
    Operation_IFC mod_445_inner <- mkRepeatStatic(8);
    Operation_IFC mod_445 <- mkDebugOperation(mod_445_inner, "mod_445");
    Operation_IFC mod_446_inner <- mkFlatten(1);
    Operation_IFC mod_446 <- mkDebugOperation(mod_446_inner, "mod_446");
    Operation_IFC mod_447_inner <- mkFlatten(0);
    Operation_IFC mod_447 <- mkDebugOperation(mod_447_inner, "mod_447");
    Operation_IFC mod_448_inner <- mkRepeatStatic(16);
    Operation_IFC mod_448 <- mkDebugOperation(mod_448_inner, "mod_448");
    Operation_IFC mod_449_inner <- mkRepeatStatic(2);
    Operation_IFC mod_449 <- mkDebugOperation(mod_449_inner, "mod_449");
    PMU_IFC mod_450_bufferize <- mkPMU(2);
    Operation_IFC mod_450_inner = mod_450_bufferize.operation;
    Operation_IFC mod_450 <- mkDebugOperation(mod_450_inner, "mod_450");
    rule rule_531;
        ChannelMessage t;
        t <- mod_433.get(0);
        mod_432.put(0, t);
    endrule
    rule rule_532;
        ChannelMessage t;
        t <- mod_416.get(1);
        mod_417.put(0, t);
    endrule
    rule rule_533;
        ChannelMessage t;
        t <- mod_414.get(1);
        mod_415.put(0, t);
    endrule
    rule rule_534;
        ChannelMessage t;
        t <- mod_426.get(1);
        mod_427.put(1, t);
    endrule
    rule rule_535;
        ChannelMessage t;
        t <- mod_432.get(0);
        mod_430.put(0, t);
    endrule
    rule rule_536;
        ChannelMessage t;
        t <- mod_442.get(1);
        mod_437.put(0, t);
    endrule
    rule rule_537;
        ChannelMessage t;
        t <- mod_444.get(0);
        mod_445.put(0, t);
    endrule
    rule rule_538;
        ChannelMessage t;
        t <- mod_450.get(1);
        mod_414.put(1, t);
    endrule
    rule rule_539;
        ChannelMessage t;
        t <- mod_428.get(1);
        mod_426.put(1, t);
    endrule
    rule rule_540;
        ChannelMessage t;
        t <- mod_431.get(0);
        mod_430.put(1, t);
    endrule
    rule rule_541;
        ChannelMessage t;
        t <- mod_436.get(0);
        mod_435.put(0, t);
    endrule
    rule rule_542;
        ChannelMessage t;
        t <- mod_420.get(0);
        mod_421.put(0, t);
    endrule
    rule rule_543;
        ChannelMessage t;
        t <- mod_412.get(0);
        mod_413.put(0, t);
    endrule
    rule rule_544;
        ChannelMessage t;
        t <- mod_430.get(0);
        mod_431.put(0, t);
    endrule
    rule rule_545;
        ChannelMessage t;
        t <- mod_440.get(0);
        mod_438.put(0, t);
    endrule
    rule rule_546;
        ChannelMessage t;
        t <- mod_435.get(0);
        mod_421.put(1, t);
    endrule
    rule rule_547;
        ChannelMessage t;
        t <- mod_422.get(0);
        mod_434.put(0, t);
    endrule
    rule rule_548;
        ChannelMessage t;
        t <- mod_421.get(0);
        mod_422.put(0, t);
    endrule
    rule rule_549;
        ChannelMessage t;
        t <- mod_425.get(0);
        mod_429.put(0, t);
    endrule
    rule rule_550;
        ChannelMessage t;
        t <- mod_448.get(0);
        mod_418.put(1, t);
    endrule
    rule rule_551;
        ChannelMessage t;
        t <- mod_416.get(0);
        mod_449.put(0, t);
    endrule
    rule rule_552;
        ChannelMessage t;
        t <- mod_449.get(0);
        mod_416.put(1, t);
    endrule
    rule rule_553;
        ChannelMessage t;
        t <- mod_434.get(0);
        mod_422.put(1, t);
    endrule
    rule rule_554;
        ChannelMessage t;
        t <- mod_447.get(0);
        mod_446.put(0, t);
    endrule
    rule rule_555;
        ChannelMessage t;
        t <- mod_438.get(0);
        mod_439.put(0, t);
    endrule
    rule rule_556;
        ChannelMessage t;
        t <- mod_438.get(1);
        mod_437.put(1, t);
    endrule
    rule rule_557;
        ChannelMessage t;
        t <- mod_443.get(0);
        mod_442.put(1, t);
    endrule
    rule rule_558;
        ChannelMessage t;
        t <- mod_417.get(1);
        mod_418.put(0, t);
    endrule
    rule rule_559;
        ChannelMessage t;
        t <- mod_418.get(1);
        mod_419.put(0, t);
    endrule
    rule rule_560;
        ChannelMessage t;
        t <- mod_417.get(0);
        mod_442.put(0, t);
    endrule
    rule rule_561;
        ChannelMessage t;
        t <- mod_419.get(0);
        mod_420.put(0, t);
    endrule
    rule rule_562;
        ChannelMessage t;
        t <- mod_430.get(1);
        mod_423.put(1, t);
    endrule
    rule rule_563;
        ChannelMessage t;
        t <- mod_425.get(1);
        mod_426.put(0, t);
    endrule
    rule rule_564;
        ChannelMessage t;
        t <- mod_429.get(0);
        mod_429.put(1, t);
    endrule
    rule rule_565;
        ChannelMessage t;
        t <- mod_437.get(0);
        mod_436.put(0, t);
    endrule
    rule rule_566;
        ChannelMessage t;
        t <- mod_439.get(0);
        mod_438.put(1, t);
    endrule
    rule rule_567;
        ChannelMessage t;
        t <- mod_442.get(0);
        mod_443.put(0, t);
    endrule
    rule rule_568;
        ChannelMessage t;
        t <- mod_422.get(1);
        mod_423.put(0, t);
    endrule
    rule rule_569;
        ChannelMessage t;
        t <- mod_414.get(0);
        mod_450.put(0, t);
    endrule
    rule rule_570;
        ChannelMessage t;
        t <- mod_411.get(0);
        mod_412.put(0, t);
    endrule
    rule rule_571;
        ChannelMessage t;
        t <- mod_415.get(3);
        mod_416.put(0, t);
    endrule
    rule rule_572;
        ChannelMessage t;
        t <- mod_413.get(0);
        mod_414.put(0, t);
    endrule
    rule rule_573;
        ChannelMessage t;
        t <- mod_441.get(0);
        mod_440.put(0, t);
    endrule
    rule rule_574;
        ChannelMessage t;
        t <- mod_446.get(0);
        mod_444.put(0, t);
    endrule
    rule rule_575;
        ChannelMessage t;
        t <- mod_429.get(1);
        mod_425.put(1, t);
    endrule
    rule rule_576;
        ChannelMessage t;
        t <- mod_426.get(0);
        mod_428.put(0, t);
    endrule
    rule rule_577;
        ChannelMessage t;
        t <- mod_418.get(0);
        mod_448.put(0, t);
    endrule
    rule rule_578;
        ChannelMessage t;
        t <- mod_444.get(1);
        mod_419.put(1, t);
    endrule
    rule rule_579;
        ChannelMessage t;
        t <- mod_450.get(0);
        mod_450.put(1, t);
    endrule
    rule rule_580;
        ChannelMessage t;
        t <- mod_424.get(0);
        mod_425.put(0, t);
    endrule
    rule rule_581;
        ChannelMessage t;
        t <- mod_423.get(0);
        mod_424.put(0, t);
    endrule
    rule rule_582;
        ChannelMessage t;
        t <- mod_445.get(0);
        mod_444.put(1, t);
    endrule
    rule rule_583;
        ChannelMessage t;
        t <- mod_428.get(0);
        mod_428.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_411.put(0, t);
        end
        if (i == 1) begin
            mod_427.put(0, t);
        end
        if (i == 2) begin
            mod_433.put(0, t);
        end
        if (i == 3) begin
            mod_441.put(0, t);
        end
        if (i == 4) begin
            mod_447.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_415.get(0);
        end
        if (i == 0) begin
            t <- mod_415.get(1);
        end
        if (i == 3) begin
            t <- mod_415.get(2);
        end
        if (i == 2) begin
            t <- mod_427.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6045 (Operation_IFC);
    Operation_IFC mod_452_inner <- mkReshape(2, 64);
    Operation_IFC mod_452 <- mkDebugOperation(mod_452_inner, "mod_452");
    Operation_IFC mod_453_inner <- mkFlatten(1);
    Operation_IFC mod_453 <- mkDebugOperation(mod_453_inner, "mod_453");
    Operation_IFC mod_454_inner <- mkFlatten(2);
    Operation_IFC mod_454 <- mkDebugOperation(mod_454_inner, "mod_454");
    Operation_IFC mod_455_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_455 <- mkDebugOperation(mod_455_inner, "mod_455");
    Broadcast_IFC#(4) mod_456_inner <- mkBroadcast(4);
    Operation_IFC mod_456 <- mkDebugOperation(mod_456_inner.op, "mod_456");
    PMU_IFC mod_457_bufferize <- mkPMU(2);
    Operation_IFC mod_457_inner = mod_457_bufferize.operation;
    Operation_IFC mod_457 <- mkDebugOperation(mod_457_inner, "mod_457");
    Broadcast_IFC#(2) mod_458_inner <- mkBroadcast(2);
    Operation_IFC mod_458 <- mkDebugOperation(mod_458_inner.op, "mod_458");
    PMU_IFC mod_459_bufferize <- mkPMU(1);
    Operation_IFC mod_459_inner = mod_459_bufferize.operation;
    Operation_IFC mod_459 <- mkDebugOperation(mod_459_inner, "mod_459");
    Operation_IFC mod_460_inner <- mkBinaryMap(1145, matmul_t_tile);
    Operation_IFC mod_460 <- mkDebugOperation(mod_460_inner, "mod_460");
    Operation_IFC mod_461_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_461 <- mkDebugOperation(mod_461_inner, "mod_461");
    Operation_IFC mod_462_inner <- mkBinaryMap(1913, mul_tile);
    Operation_IFC mod_462 <- mkDebugOperation(mod_462_inner, "mod_462");
    PMU_IFC mod_463_bufferize <- mkPMU(1);
    Operation_IFC mod_463_inner = mod_463_bufferize.operation;
    Operation_IFC mod_463 <- mkDebugOperation(mod_463_inner, "mod_463");
    Operation_IFC mod_464_inner <- mkBinaryMap(2541, matmul_t_tile);
    Operation_IFC mod_464 <- mkDebugOperation(mod_464_inner, "mod_464");
    Operation_IFC mod_465_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_465 <- mkDebugOperation(mod_465_inner, "mod_465");
    Operation_IFC mod_466_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_466 <- mkDebugOperation(mod_466_inner, "mod_466");
    Operation_IFC mod_467_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_467 <- mkDebugOperation(mod_467_inner, "mod_467");
    Operation_IFC mod_468_inner <- mkBinaryMap(2812, mul_tile);
    Operation_IFC mod_468 <- mkDebugOperation(mod_468_inner, "mod_468");
    PMU_IFC mod_469_bufferize <- mkPMU(1);
    Operation_IFC mod_469_inner = mod_469_bufferize.operation;
    Operation_IFC mod_469 <- mkDebugOperation(mod_469_inner, "mod_469");
    PMU_IFC mod_470_bufferize <- mkPMU(2);
    Operation_IFC mod_470_inner = mod_470_bufferize.operation;
    Operation_IFC mod_470 <- mkDebugOperation(mod_470_inner, "mod_470");
    PMU_IFC mod_471_bufferize <- mkPMU(2);
    Operation_IFC mod_471_inner = mod_471_bufferize.operation;
    Operation_IFC mod_471 <- mkDebugOperation(mod_471_inner, "mod_471");
    Operation_IFC mod_472_inner <- mkRepeatStatic(8);
    Operation_IFC mod_472 <- mkDebugOperation(mod_472_inner, "mod_472");
    Operation_IFC mod_473_inner <- mkFlatten(1);
    Operation_IFC mod_473 <- mkDebugOperation(mod_473_inner, "mod_473");
    Operation_IFC mod_474_inner <- mkFlatten(0);
    Operation_IFC mod_474 <- mkDebugOperation(mod_474_inner, "mod_474");
    Operation_IFC mod_475_inner <- mkRepeatStatic(3);
    Operation_IFC mod_475 <- mkDebugOperation(mod_475_inner, "mod_475");
    Operation_IFC mod_476_inner <- mkUnaryMap(1785, silu_tile);
    Operation_IFC mod_476 <- mkDebugOperation(mod_476_inner, "mod_476");
    Operation_IFC mod_477_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_477 <- mkDebugOperation(mod_477_inner, "mod_477");
    Operation_IFC mod_478_inner <- mkBinaryMap(1657, matmul_t_tile);
    Operation_IFC mod_478 <- mkDebugOperation(mod_478_inner, "mod_478");
    PMU_IFC mod_479_bufferize <- mkPMU(2);
    Operation_IFC mod_479_inner = mod_479_bufferize.operation;
    Operation_IFC mod_479 <- mkDebugOperation(mod_479_inner, "mod_479");
    Operation_IFC mod_480_inner <- mkRepeatStatic(8);
    Operation_IFC mod_480 <- mkDebugOperation(mod_480_inner, "mod_480");
    Operation_IFC mod_481_inner <- mkFlatten(1);
    Operation_IFC mod_481 <- mkDebugOperation(mod_481_inner, "mod_481");
    Operation_IFC mod_482_inner <- mkFlatten(0);
    Operation_IFC mod_482 <- mkDebugOperation(mod_482_inner, "mod_482");
    PMU_IFC mod_483_bufferize <- mkPMU(1);
    Operation_IFC mod_483_inner = mod_483_bufferize.operation;
    Operation_IFC mod_483 <- mkDebugOperation(mod_483_inner, "mod_483");
    Operation_IFC mod_484_inner <- mkRepeatStatic(16);
    Operation_IFC mod_484 <- mkDebugOperation(mod_484_inner, "mod_484");
    PMU_IFC mod_485_bufferize <- mkPMU(2);
    Operation_IFC mod_485_inner = mod_485_bufferize.operation;
    Operation_IFC mod_485 <- mkDebugOperation(mod_485_inner, "mod_485");
    Operation_IFC mod_486_inner <- mkRepeatStatic(8);
    Operation_IFC mod_486 <- mkDebugOperation(mod_486_inner, "mod_486");
    Operation_IFC mod_487_inner <- mkFlatten(1);
    Operation_IFC mod_487 <- mkDebugOperation(mod_487_inner, "mod_487");
    Operation_IFC mod_488_inner <- mkFlatten(0);
    Operation_IFC mod_488 <- mkDebugOperation(mod_488_inner, "mod_488");
    Operation_IFC mod_489_inner <- mkRepeatStatic(16);
    Operation_IFC mod_489 <- mkDebugOperation(mod_489_inner, "mod_489");
    Operation_IFC mod_490_inner <- mkRepeatStatic(2);
    Operation_IFC mod_490 <- mkDebugOperation(mod_490_inner, "mod_490");
    PMU_IFC mod_491_bufferize <- mkPMU(2);
    Operation_IFC mod_491_inner = mod_491_bufferize.operation;
    Operation_IFC mod_491 <- mkDebugOperation(mod_491_inner, "mod_491");
    rule rule_584;
        ChannelMessage t;
        t <- mod_490.get(0);
        mod_457.put(1, t);
    endrule
    rule rule_585;
        ChannelMessage t;
        t <- mod_474.get(0);
        mod_473.put(0, t);
    endrule
    rule rule_586;
        ChannelMessage t;
        t <- mod_471.get(1);
        mod_464.put(1, t);
    endrule
    rule rule_587;
        ChannelMessage t;
        t <- mod_466.get(1);
        mod_467.put(0, t);
    endrule
    rule rule_588;
        ChannelMessage t;
        t <- mod_484.get(0);
        mod_483.put(1, t);
    endrule
    rule rule_589;
        ChannelMessage t;
        t <- mod_463.get(1);
        mod_464.put(0, t);
    endrule
    rule rule_590;
        ChannelMessage t;
        t <- mod_457.get(1);
        mod_458.put(0, t);
    endrule
    rule rule_591;
        ChannelMessage t;
        t <- mod_483.get(1);
        mod_478.put(0, t);
    endrule
    rule rule_592;
        ChannelMessage t;
        t <- mod_455.get(1);
        mod_456.put(0, t);
    endrule
    rule rule_593;
        ChannelMessage t;
        t <- mod_485.get(1);
        mod_460.put(1, t);
    endrule
    rule rule_594;
        ChannelMessage t;
        t <- mod_457.get(0);
        mod_490.put(0, t);
    endrule
    rule rule_595;
        ChannelMessage t;
        t <- mod_466.get(0);
        mod_470.put(0, t);
    endrule
    rule rule_596;
        ChannelMessage t;
        t <- mod_455.get(0);
        mod_491.put(0, t);
    endrule
    rule rule_597;
        ChannelMessage t;
        t <- mod_480.get(0);
        mod_479.put(1, t);
    endrule
    rule rule_598;
        ChannelMessage t;
        t <- mod_472.get(0);
        mod_471.put(1, t);
    endrule
    rule rule_599;
        ChannelMessage t;
        t <- mod_483.get(0);
        mod_484.put(0, t);
    endrule
    rule rule_600;
        ChannelMessage t;
        t <- mod_489.get(0);
        mod_459.put(1, t);
    endrule
    rule rule_601;
        ChannelMessage t;
        t <- mod_491.get(0);
        mod_491.put(1, t);
    endrule
    rule rule_602;
        ChannelMessage t;
        t <- mod_491.get(1);
        mod_455.put(1, t);
    endrule
    rule rule_603;
        ChannelMessage t;
        t <- mod_465.get(0);
        mod_466.put(0, t);
    endrule
    rule rule_604;
        ChannelMessage t;
        t <- mod_454.get(0);
        mod_455.put(0, t);
    endrule
    rule rule_605;
        ChannelMessage t;
        t <- mod_453.get(0);
        mod_454.put(0, t);
    endrule
    rule rule_606;
        ChannelMessage t;
        t <- mod_469.get(0);
        mod_469.put(1, t);
    endrule
    rule rule_607;
        ChannelMessage t;
        t <- mod_471.get(0);
        mod_472.put(0, t);
    endrule
    rule rule_608;
        ChannelMessage t;
        t <- mod_467.get(1);
        mod_468.put(1, t);
    endrule
    rule rule_609;
        ChannelMessage t;
        t <- mod_476.get(0);
        mod_462.put(1, t);
    endrule
    rule rule_610;
        ChannelMessage t;
        t <- mod_458.get(0);
        mod_483.put(0, t);
    endrule
    rule rule_611;
        ChannelMessage t;
        t <- mod_459.get(0);
        mod_489.put(0, t);
    endrule
    rule rule_612;
        ChannelMessage t;
        t <- mod_470.get(0);
        mod_470.put(1, t);
    endrule
    rule rule_613;
        ChannelMessage t;
        t <- mod_464.get(0);
        mod_465.put(0, t);
    endrule
    rule rule_614;
        ChannelMessage t;
        t <- mod_475.get(0);
        mod_463.put(1, t);
    endrule
    rule rule_615;
        ChannelMessage t;
        t <- mod_459.get(1);
        mod_460.put(0, t);
    endrule
    rule rule_616;
        ChannelMessage t;
        t <- mod_461.get(0);
        mod_462.put(0, t);
    endrule
    rule rule_617;
        ChannelMessage t;
        t <- mod_460.get(0);
        mod_461.put(0, t);
    endrule
    rule rule_618;
        ChannelMessage t;
        t <- mod_481.get(0);
        mod_479.put(0, t);
    endrule
    rule rule_619;
        ChannelMessage t;
        t <- mod_473.get(0);
        mod_471.put(0, t);
    endrule
    rule rule_620;
        ChannelMessage t;
        t <- mod_462.get(0);
        mod_463.put(0, t);
    endrule
    rule rule_621;
        ChannelMessage t;
        t <- mod_482.get(0);
        mod_481.put(0, t);
    endrule
    rule rule_622;
        ChannelMessage t;
        t <- mod_486.get(0);
        mod_485.put(1, t);
    endrule
    rule rule_623;
        ChannelMessage t;
        t <- mod_488.get(0);
        mod_487.put(0, t);
    endrule
    rule rule_624;
        ChannelMessage t;
        t <- mod_479.get(0);
        mod_480.put(0, t);
    endrule
    rule rule_625;
        ChannelMessage t;
        t <- mod_458.get(1);
        mod_459.put(0, t);
    endrule
    rule rule_626;
        ChannelMessage t;
        t <- mod_467.get(0);
        mod_469.put(0, t);
    endrule
    rule rule_627;
        ChannelMessage t;
        t <- mod_470.get(1);
        mod_466.put(1, t);
    endrule
    rule rule_628;
        ChannelMessage t;
        t <- mod_452.get(0);
        mod_453.put(0, t);
    endrule
    rule rule_629;
        ChannelMessage t;
        t <- mod_469.get(1);
        mod_467.put(1, t);
    endrule
    rule rule_630;
        ChannelMessage t;
        t <- mod_487.get(0);
        mod_485.put(0, t);
    endrule
    rule rule_631;
        ChannelMessage t;
        t <- mod_463.get(0);
        mod_475.put(0, t);
    endrule
    rule rule_632;
        ChannelMessage t;
        t <- mod_456.get(3);
        mod_457.put(0, t);
    endrule
    rule rule_633;
        ChannelMessage t;
        t <- mod_485.get(0);
        mod_486.put(0, t);
    endrule
    rule rule_634;
        ChannelMessage t;
        t <- mod_478.get(0);
        mod_477.put(0, t);
    endrule
    rule rule_635;
        ChannelMessage t;
        t <- mod_479.get(1);
        mod_478.put(1, t);
    endrule
    rule rule_636;
        ChannelMessage t;
        t <- mod_477.get(0);
        mod_476.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_452.put(0, t);
        end
        if (i == 1) begin
            mod_468.put(0, t);
        end
        if (i == 2) begin
            mod_474.put(0, t);
        end
        if (i == 3) begin
            mod_482.put(0, t);
        end
        if (i == 4) begin
            mod_488.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_456.get(0);
        end
        if (i == 0) begin
            t <- mod_456.get(1);
        end
        if (i == 2) begin
            t <- mod_456.get(2);
        end
        if (i == 1) begin
            t <- mod_468.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6046 (Operation_IFC);
    Operation_IFC mod_493_inner <- mkReshape(2, 64);
    Operation_IFC mod_493 <- mkDebugOperation(mod_493_inner, "mod_493");
    Operation_IFC mod_494_inner <- mkFlatten(1);
    Operation_IFC mod_494 <- mkDebugOperation(mod_494_inner, "mod_494");
    Operation_IFC mod_495_inner <- mkFlatten(2);
    Operation_IFC mod_495 <- mkDebugOperation(mod_495_inner, "mod_495");
    Operation_IFC mod_496_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_496 <- mkDebugOperation(mod_496_inner, "mod_496");
    Broadcast_IFC#(4) mod_497_inner <- mkBroadcast(4);
    Operation_IFC mod_497 <- mkDebugOperation(mod_497_inner.op, "mod_497");
    PMU_IFC mod_498_bufferize <- mkPMU(2);
    Operation_IFC mod_498_inner = mod_498_bufferize.operation;
    Operation_IFC mod_498 <- mkDebugOperation(mod_498_inner, "mod_498");
    Broadcast_IFC#(2) mod_499_inner <- mkBroadcast(2);
    Operation_IFC mod_499 <- mkDebugOperation(mod_499_inner.op, "mod_499");
    PMU_IFC mod_500_bufferize <- mkPMU(1);
    Operation_IFC mod_500_inner = mod_500_bufferize.operation;
    Operation_IFC mod_500 <- mkDebugOperation(mod_500_inner, "mod_500");
    Operation_IFC mod_501_inner <- mkBinaryMap(1144, matmul_t_tile);
    Operation_IFC mod_501 <- mkDebugOperation(mod_501_inner, "mod_501");
    Operation_IFC mod_502_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_502 <- mkDebugOperation(mod_502_inner, "mod_502");
    Operation_IFC mod_503_inner <- mkBinaryMap(1912, mul_tile);
    Operation_IFC mod_503 <- mkDebugOperation(mod_503_inner, "mod_503");
    PMU_IFC mod_504_bufferize <- mkPMU(1);
    Operation_IFC mod_504_inner = mod_504_bufferize.operation;
    Operation_IFC mod_504 <- mkDebugOperation(mod_504_inner, "mod_504");
    Operation_IFC mod_505_inner <- mkBinaryMap(2539, matmul_t_tile);
    Operation_IFC mod_505 <- mkDebugOperation(mod_505_inner, "mod_505");
    Operation_IFC mod_506_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_506 <- mkDebugOperation(mod_506_inner, "mod_506");
    Operation_IFC mod_507_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_507 <- mkDebugOperation(mod_507_inner, "mod_507");
    Operation_IFC mod_508_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_508 <- mkDebugOperation(mod_508_inner, "mod_508");
    Operation_IFC mod_509_inner <- mkBinaryMap(2811, mul_tile);
    Operation_IFC mod_509 <- mkDebugOperation(mod_509_inner, "mod_509");
    PMU_IFC mod_510_bufferize <- mkPMU(1);
    Operation_IFC mod_510_inner = mod_510_bufferize.operation;
    Operation_IFC mod_510 <- mkDebugOperation(mod_510_inner, "mod_510");
    PMU_IFC mod_511_bufferize <- mkPMU(2);
    Operation_IFC mod_511_inner = mod_511_bufferize.operation;
    Operation_IFC mod_511 <- mkDebugOperation(mod_511_inner, "mod_511");
    PMU_IFC mod_512_bufferize <- mkPMU(2);
    Operation_IFC mod_512_inner = mod_512_bufferize.operation;
    Operation_IFC mod_512 <- mkDebugOperation(mod_512_inner, "mod_512");
    Operation_IFC mod_513_inner <- mkRepeatStatic(8);
    Operation_IFC mod_513 <- mkDebugOperation(mod_513_inner, "mod_513");
    Operation_IFC mod_514_inner <- mkFlatten(1);
    Operation_IFC mod_514 <- mkDebugOperation(mod_514_inner, "mod_514");
    Operation_IFC mod_515_inner <- mkFlatten(0);
    Operation_IFC mod_515 <- mkDebugOperation(mod_515_inner, "mod_515");
    Operation_IFC mod_516_inner <- mkRepeatStatic(3);
    Operation_IFC mod_516 <- mkDebugOperation(mod_516_inner, "mod_516");
    Operation_IFC mod_517_inner <- mkUnaryMap(1784, silu_tile);
    Operation_IFC mod_517 <- mkDebugOperation(mod_517_inner, "mod_517");
    Operation_IFC mod_518_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_518 <- mkDebugOperation(mod_518_inner, "mod_518");
    Operation_IFC mod_519_inner <- mkBinaryMap(1656, matmul_t_tile);
    Operation_IFC mod_519 <- mkDebugOperation(mod_519_inner, "mod_519");
    PMU_IFC mod_520_bufferize <- mkPMU(2);
    Operation_IFC mod_520_inner = mod_520_bufferize.operation;
    Operation_IFC mod_520 <- mkDebugOperation(mod_520_inner, "mod_520");
    Operation_IFC mod_521_inner <- mkRepeatStatic(8);
    Operation_IFC mod_521 <- mkDebugOperation(mod_521_inner, "mod_521");
    Operation_IFC mod_522_inner <- mkFlatten(1);
    Operation_IFC mod_522 <- mkDebugOperation(mod_522_inner, "mod_522");
    Operation_IFC mod_523_inner <- mkFlatten(0);
    Operation_IFC mod_523 <- mkDebugOperation(mod_523_inner, "mod_523");
    PMU_IFC mod_524_bufferize <- mkPMU(1);
    Operation_IFC mod_524_inner = mod_524_bufferize.operation;
    Operation_IFC mod_524 <- mkDebugOperation(mod_524_inner, "mod_524");
    Operation_IFC mod_525_inner <- mkRepeatStatic(16);
    Operation_IFC mod_525 <- mkDebugOperation(mod_525_inner, "mod_525");
    PMU_IFC mod_526_bufferize <- mkPMU(2);
    Operation_IFC mod_526_inner = mod_526_bufferize.operation;
    Operation_IFC mod_526 <- mkDebugOperation(mod_526_inner, "mod_526");
    Operation_IFC mod_527_inner <- mkRepeatStatic(8);
    Operation_IFC mod_527 <- mkDebugOperation(mod_527_inner, "mod_527");
    Operation_IFC mod_528_inner <- mkFlatten(1);
    Operation_IFC mod_528 <- mkDebugOperation(mod_528_inner, "mod_528");
    Operation_IFC mod_529_inner <- mkFlatten(0);
    Operation_IFC mod_529 <- mkDebugOperation(mod_529_inner, "mod_529");
    Operation_IFC mod_530_inner <- mkRepeatStatic(16);
    Operation_IFC mod_530 <- mkDebugOperation(mod_530_inner, "mod_530");
    Operation_IFC mod_531_inner <- mkRepeatStatic(2);
    Operation_IFC mod_531 <- mkDebugOperation(mod_531_inner, "mod_531");
    PMU_IFC mod_532_bufferize <- mkPMU(2);
    Operation_IFC mod_532_inner = mod_532_bufferize.operation;
    Operation_IFC mod_532 <- mkDebugOperation(mod_532_inner, "mod_532");
    rule rule_637;
        ChannelMessage t;
        t <- mod_513.get(0);
        mod_512.put(1, t);
    endrule
    rule rule_638;
        ChannelMessage t;
        t <- mod_510.get(0);
        mod_510.put(1, t);
    endrule
    rule rule_639;
        ChannelMessage t;
        t <- mod_494.get(0);
        mod_495.put(0, t);
    endrule
    rule rule_640;
        ChannelMessage t;
        t <- mod_498.get(1);
        mod_499.put(0, t);
    endrule
    rule rule_641;
        ChannelMessage t;
        t <- mod_520.get(0);
        mod_521.put(0, t);
    endrule
    rule rule_642;
        ChannelMessage t;
        t <- mod_500.get(1);
        mod_501.put(0, t);
    endrule
    rule rule_643;
        ChannelMessage t;
        t <- mod_496.get(1);
        mod_497.put(0, t);
    endrule
    rule rule_644;
        ChannelMessage t;
        t <- mod_508.get(0);
        mod_510.put(0, t);
    endrule
    rule rule_645;
        ChannelMessage t;
        t <- mod_511.get(1);
        mod_507.put(1, t);
    endrule
    rule rule_646;
        ChannelMessage t;
        t <- mod_514.get(0);
        mod_512.put(0, t);
    endrule
    rule rule_647;
        ChannelMessage t;
        t <- mod_506.get(0);
        mod_507.put(0, t);
    endrule
    rule rule_648;
        ChannelMessage t;
        t <- mod_501.get(0);
        mod_502.put(0, t);
    endrule
    rule rule_649;
        ChannelMessage t;
        t <- mod_525.get(0);
        mod_524.put(1, t);
    endrule
    rule rule_650;
        ChannelMessage t;
        t <- mod_532.get(0);
        mod_532.put(1, t);
    endrule
    rule rule_651;
        ChannelMessage t;
        t <- mod_531.get(0);
        mod_498.put(1, t);
    endrule
    rule rule_652;
        ChannelMessage t;
        t <- mod_517.get(0);
        mod_503.put(1, t);
    endrule
    rule rule_653;
        ChannelMessage t;
        t <- mod_493.get(0);
        mod_494.put(0, t);
    endrule
    rule rule_654;
        ChannelMessage t;
        t <- mod_498.get(0);
        mod_531.put(0, t);
    endrule
    rule rule_655;
        ChannelMessage t;
        t <- mod_510.get(1);
        mod_508.put(1, t);
    endrule
    rule rule_656;
        ChannelMessage t;
        t <- mod_504.get(1);
        mod_505.put(0, t);
    endrule
    rule rule_657;
        ChannelMessage t;
        t <- mod_507.get(1);
        mod_508.put(0, t);
    endrule
    rule rule_658;
        ChannelMessage t;
        t <- mod_497.get(3);
        mod_498.put(0, t);
    endrule
    rule rule_659;
        ChannelMessage t;
        t <- mod_499.get(0);
        mod_524.put(0, t);
    endrule
    rule rule_660;
        ChannelMessage t;
        t <- mod_521.get(0);
        mod_520.put(1, t);
    endrule
    rule rule_661;
        ChannelMessage t;
        t <- mod_529.get(0);
        mod_528.put(0, t);
    endrule
    rule rule_662;
        ChannelMessage t;
        t <- mod_520.get(1);
        mod_519.put(1, t);
    endrule
    rule rule_663;
        ChannelMessage t;
        t <- mod_526.get(0);
        mod_527.put(0, t);
    endrule
    rule rule_664;
        ChannelMessage t;
        t <- mod_526.get(1);
        mod_501.put(1, t);
    endrule
    rule rule_665;
        ChannelMessage t;
        t <- mod_508.get(1);
        mod_509.put(1, t);
    endrule
    rule rule_666;
        ChannelMessage t;
        t <- mod_522.get(0);
        mod_520.put(0, t);
    endrule
    rule rule_667;
        ChannelMessage t;
        t <- mod_499.get(1);
        mod_500.put(0, t);
    endrule
    rule rule_668;
        ChannelMessage t;
        t <- mod_512.get(1);
        mod_505.put(1, t);
    endrule
    rule rule_669;
        ChannelMessage t;
        t <- mod_530.get(0);
        mod_500.put(1, t);
    endrule
    rule rule_670;
        ChannelMessage t;
        t <- mod_495.get(0);
        mod_496.put(0, t);
    endrule
    rule rule_671;
        ChannelMessage t;
        t <- mod_502.get(0);
        mod_503.put(0, t);
    endrule
    rule rule_672;
        ChannelMessage t;
        t <- mod_505.get(0);
        mod_506.put(0, t);
    endrule
    rule rule_673;
        ChannelMessage t;
        t <- mod_523.get(0);
        mod_522.put(0, t);
    endrule
    rule rule_674;
        ChannelMessage t;
        t <- mod_511.get(0);
        mod_511.put(1, t);
    endrule
    rule rule_675;
        ChannelMessage t;
        t <- mod_524.get(1);
        mod_519.put(0, t);
    endrule
    rule rule_676;
        ChannelMessage t;
        t <- mod_515.get(0);
        mod_514.put(0, t);
    endrule
    rule rule_677;
        ChannelMessage t;
        t <- mod_519.get(0);
        mod_518.put(0, t);
    endrule
    rule rule_678;
        ChannelMessage t;
        t <- mod_532.get(1);
        mod_496.put(1, t);
    endrule
    rule rule_679;
        ChannelMessage t;
        t <- mod_516.get(0);
        mod_504.put(1, t);
    endrule
    rule rule_680;
        ChannelMessage t;
        t <- mod_512.get(0);
        mod_513.put(0, t);
    endrule
    rule rule_681;
        ChannelMessage t;
        t <- mod_500.get(0);
        mod_530.put(0, t);
    endrule
    rule rule_682;
        ChannelMessage t;
        t <- mod_518.get(0);
        mod_517.put(0, t);
    endrule
    rule rule_683;
        ChannelMessage t;
        t <- mod_503.get(0);
        mod_504.put(0, t);
    endrule
    rule rule_684;
        ChannelMessage t;
        t <- mod_507.get(0);
        mod_511.put(0, t);
    endrule
    rule rule_685;
        ChannelMessage t;
        t <- mod_524.get(0);
        mod_525.put(0, t);
    endrule
    rule rule_686;
        ChannelMessage t;
        t <- mod_504.get(0);
        mod_516.put(0, t);
    endrule
    rule rule_687;
        ChannelMessage t;
        t <- mod_496.get(0);
        mod_532.put(0, t);
    endrule
    rule rule_688;
        ChannelMessage t;
        t <- mod_527.get(0);
        mod_526.put(1, t);
    endrule
    rule rule_689;
        ChannelMessage t;
        t <- mod_528.get(0);
        mod_526.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_493.put(0, t);
        end
        if (i == 1) begin
            mod_509.put(0, t);
        end
        if (i == 2) begin
            mod_515.put(0, t);
        end
        if (i == 3) begin
            mod_523.put(0, t);
        end
        if (i == 4) begin
            mod_529.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_497.get(0);
        end
        if (i == 2) begin
            t <- mod_497.get(1);
        end
        if (i == 3) begin
            t <- mod_497.get(2);
        end
        if (i == 1) begin
            t <- mod_509.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6047 (Operation_IFC);
    Operation_IFC mod_534_inner <- mkReshape(2, 64);
    Operation_IFC mod_534 <- mkDebugOperation(mod_534_inner, "mod_534");
    Operation_IFC mod_535_inner <- mkFlatten(1);
    Operation_IFC mod_535 <- mkDebugOperation(mod_535_inner, "mod_535");
    Operation_IFC mod_536_inner <- mkFlatten(2);
    Operation_IFC mod_536 <- mkDebugOperation(mod_536_inner, "mod_536");
    Operation_IFC mod_537_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_537 <- mkDebugOperation(mod_537_inner, "mod_537");
    Broadcast_IFC#(4) mod_538_inner <- mkBroadcast(4);
    Operation_IFC mod_538 <- mkDebugOperation(mod_538_inner.op, "mod_538");
    PMU_IFC mod_539_bufferize <- mkPMU(2);
    Operation_IFC mod_539_inner = mod_539_bufferize.operation;
    Operation_IFC mod_539 <- mkDebugOperation(mod_539_inner, "mod_539");
    Broadcast_IFC#(2) mod_540_inner <- mkBroadcast(2);
    Operation_IFC mod_540 <- mkDebugOperation(mod_540_inner.op, "mod_540");
    PMU_IFC mod_541_bufferize <- mkPMU(1);
    Operation_IFC mod_541_inner = mod_541_bufferize.operation;
    Operation_IFC mod_541 <- mkDebugOperation(mod_541_inner, "mod_541");
    Operation_IFC mod_542_inner <- mkBinaryMap(1143, matmul_t_tile);
    Operation_IFC mod_542 <- mkDebugOperation(mod_542_inner, "mod_542");
    Operation_IFC mod_543_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_543 <- mkDebugOperation(mod_543_inner, "mod_543");
    Operation_IFC mod_544_inner <- mkBinaryMap(1911, mul_tile);
    Operation_IFC mod_544 <- mkDebugOperation(mod_544_inner, "mod_544");
    PMU_IFC mod_545_bufferize <- mkPMU(1);
    Operation_IFC mod_545_inner = mod_545_bufferize.operation;
    Operation_IFC mod_545 <- mkDebugOperation(mod_545_inner, "mod_545");
    Operation_IFC mod_546_inner <- mkBinaryMap(2537, matmul_t_tile);
    Operation_IFC mod_546 <- mkDebugOperation(mod_546_inner, "mod_546");
    Operation_IFC mod_547_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_547 <- mkDebugOperation(mod_547_inner, "mod_547");
    Operation_IFC mod_548_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_548 <- mkDebugOperation(mod_548_inner, "mod_548");
    Operation_IFC mod_549_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_549 <- mkDebugOperation(mod_549_inner, "mod_549");
    Operation_IFC mod_550_inner <- mkBinaryMap(2810, mul_tile);
    Operation_IFC mod_550 <- mkDebugOperation(mod_550_inner, "mod_550");
    PMU_IFC mod_551_bufferize <- mkPMU(1);
    Operation_IFC mod_551_inner = mod_551_bufferize.operation;
    Operation_IFC mod_551 <- mkDebugOperation(mod_551_inner, "mod_551");
    PMU_IFC mod_552_bufferize <- mkPMU(2);
    Operation_IFC mod_552_inner = mod_552_bufferize.operation;
    Operation_IFC mod_552 <- mkDebugOperation(mod_552_inner, "mod_552");
    PMU_IFC mod_553_bufferize <- mkPMU(2);
    Operation_IFC mod_553_inner = mod_553_bufferize.operation;
    Operation_IFC mod_553 <- mkDebugOperation(mod_553_inner, "mod_553");
    Operation_IFC mod_554_inner <- mkRepeatStatic(8);
    Operation_IFC mod_554 <- mkDebugOperation(mod_554_inner, "mod_554");
    Operation_IFC mod_555_inner <- mkFlatten(1);
    Operation_IFC mod_555 <- mkDebugOperation(mod_555_inner, "mod_555");
    Operation_IFC mod_556_inner <- mkFlatten(0);
    Operation_IFC mod_556 <- mkDebugOperation(mod_556_inner, "mod_556");
    Operation_IFC mod_557_inner <- mkRepeatStatic(3);
    Operation_IFC mod_557 <- mkDebugOperation(mod_557_inner, "mod_557");
    Operation_IFC mod_558_inner <- mkUnaryMap(1783, silu_tile);
    Operation_IFC mod_558 <- mkDebugOperation(mod_558_inner, "mod_558");
    Operation_IFC mod_559_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_559 <- mkDebugOperation(mod_559_inner, "mod_559");
    Operation_IFC mod_560_inner <- mkBinaryMap(1655, matmul_t_tile);
    Operation_IFC mod_560 <- mkDebugOperation(mod_560_inner, "mod_560");
    PMU_IFC mod_561_bufferize <- mkPMU(2);
    Operation_IFC mod_561_inner = mod_561_bufferize.operation;
    Operation_IFC mod_561 <- mkDebugOperation(mod_561_inner, "mod_561");
    Operation_IFC mod_562_inner <- mkRepeatStatic(8);
    Operation_IFC mod_562 <- mkDebugOperation(mod_562_inner, "mod_562");
    Operation_IFC mod_563_inner <- mkFlatten(1);
    Operation_IFC mod_563 <- mkDebugOperation(mod_563_inner, "mod_563");
    Operation_IFC mod_564_inner <- mkFlatten(0);
    Operation_IFC mod_564 <- mkDebugOperation(mod_564_inner, "mod_564");
    PMU_IFC mod_565_bufferize <- mkPMU(1);
    Operation_IFC mod_565_inner = mod_565_bufferize.operation;
    Operation_IFC mod_565 <- mkDebugOperation(mod_565_inner, "mod_565");
    Operation_IFC mod_566_inner <- mkRepeatStatic(16);
    Operation_IFC mod_566 <- mkDebugOperation(mod_566_inner, "mod_566");
    PMU_IFC mod_567_bufferize <- mkPMU(2);
    Operation_IFC mod_567_inner = mod_567_bufferize.operation;
    Operation_IFC mod_567 <- mkDebugOperation(mod_567_inner, "mod_567");
    Operation_IFC mod_568_inner <- mkRepeatStatic(8);
    Operation_IFC mod_568 <- mkDebugOperation(mod_568_inner, "mod_568");
    Operation_IFC mod_569_inner <- mkFlatten(1);
    Operation_IFC mod_569 <- mkDebugOperation(mod_569_inner, "mod_569");
    Operation_IFC mod_570_inner <- mkFlatten(0);
    Operation_IFC mod_570 <- mkDebugOperation(mod_570_inner, "mod_570");
    Operation_IFC mod_571_inner <- mkRepeatStatic(16);
    Operation_IFC mod_571 <- mkDebugOperation(mod_571_inner, "mod_571");
    Operation_IFC mod_572_inner <- mkRepeatStatic(2);
    Operation_IFC mod_572 <- mkDebugOperation(mod_572_inner, "mod_572");
    PMU_IFC mod_573_bufferize <- mkPMU(2);
    Operation_IFC mod_573_inner = mod_573_bufferize.operation;
    Operation_IFC mod_573 <- mkDebugOperation(mod_573_inner, "mod_573");
    rule rule_690;
        ChannelMessage t;
        t <- mod_568.get(0);
        mod_567.put(1, t);
    endrule
    rule rule_691;
        ChannelMessage t;
        t <- mod_540.get(1);
        mod_541.put(0, t);
    endrule
    rule rule_692;
        ChannelMessage t;
        t <- mod_569.get(0);
        mod_567.put(0, t);
    endrule
    rule rule_693;
        ChannelMessage t;
        t <- mod_566.get(0);
        mod_565.put(1, t);
    endrule
    rule rule_694;
        ChannelMessage t;
        t <- mod_537.get(1);
        mod_538.put(0, t);
    endrule
    rule rule_695;
        ChannelMessage t;
        t <- mod_544.get(0);
        mod_545.put(0, t);
    endrule
    rule rule_696;
        ChannelMessage t;
        t <- mod_543.get(0);
        mod_544.put(0, t);
    endrule
    rule rule_697;
        ChannelMessage t;
        t <- mod_552.get(1);
        mod_548.put(1, t);
    endrule
    rule rule_698;
        ChannelMessage t;
        t <- mod_554.get(0);
        mod_553.put(1, t);
    endrule
    rule rule_699;
        ChannelMessage t;
        t <- mod_561.get(0);
        mod_562.put(0, t);
    endrule
    rule rule_700;
        ChannelMessage t;
        t <- mod_564.get(0);
        mod_563.put(0, t);
    endrule
    rule rule_701;
        ChannelMessage t;
        t <- mod_570.get(0);
        mod_569.put(0, t);
    endrule
    rule rule_702;
        ChannelMessage t;
        t <- mod_571.get(0);
        mod_541.put(1, t);
    endrule
    rule rule_703;
        ChannelMessage t;
        t <- mod_536.get(0);
        mod_537.put(0, t);
    endrule
    rule rule_704;
        ChannelMessage t;
        t <- mod_556.get(0);
        mod_555.put(0, t);
    endrule
    rule rule_705;
        ChannelMessage t;
        t <- mod_548.get(1);
        mod_549.put(0, t);
    endrule
    rule rule_706;
        ChannelMessage t;
        t <- mod_565.get(0);
        mod_566.put(0, t);
    endrule
    rule rule_707;
        ChannelMessage t;
        t <- mod_542.get(0);
        mod_543.put(0, t);
    endrule
    rule rule_708;
        ChannelMessage t;
        t <- mod_541.get(0);
        mod_571.put(0, t);
    endrule
    rule rule_709;
        ChannelMessage t;
        t <- mod_551.get(0);
        mod_551.put(1, t);
    endrule
    rule rule_710;
        ChannelMessage t;
        t <- mod_573.get(0);
        mod_573.put(1, t);
    endrule
    rule rule_711;
        ChannelMessage t;
        t <- mod_551.get(1);
        mod_549.put(1, t);
    endrule
    rule rule_712;
        ChannelMessage t;
        t <- mod_573.get(1);
        mod_537.put(1, t);
    endrule
    rule rule_713;
        ChannelMessage t;
        t <- mod_545.get(0);
        mod_557.put(0, t);
    endrule
    rule rule_714;
        ChannelMessage t;
        t <- mod_547.get(0);
        mod_548.put(0, t);
    endrule
    rule rule_715;
        ChannelMessage t;
        t <- mod_560.get(0);
        mod_559.put(0, t);
    endrule
    rule rule_716;
        ChannelMessage t;
        t <- mod_565.get(1);
        mod_560.put(0, t);
    endrule
    rule rule_717;
        ChannelMessage t;
        t <- mod_546.get(0);
        mod_547.put(0, t);
    endrule
    rule rule_718;
        ChannelMessage t;
        t <- mod_549.get(1);
        mod_550.put(1, t);
    endrule
    rule rule_719;
        ChannelMessage t;
        t <- mod_537.get(0);
        mod_573.put(0, t);
    endrule
    rule rule_720;
        ChannelMessage t;
        t <- mod_540.get(0);
        mod_565.put(0, t);
    endrule
    rule rule_721;
        ChannelMessage t;
        t <- mod_558.get(0);
        mod_544.put(1, t);
    endrule
    rule rule_722;
        ChannelMessage t;
        t <- mod_559.get(0);
        mod_558.put(0, t);
    endrule
    rule rule_723;
        ChannelMessage t;
        t <- mod_572.get(0);
        mod_539.put(1, t);
    endrule
    rule rule_724;
        ChannelMessage t;
        t <- mod_534.get(0);
        mod_535.put(0, t);
    endrule
    rule rule_725;
        ChannelMessage t;
        t <- mod_553.get(0);
        mod_554.put(0, t);
    endrule
    rule rule_726;
        ChannelMessage t;
        t <- mod_539.get(1);
        mod_540.put(0, t);
    endrule
    rule rule_727;
        ChannelMessage t;
        t <- mod_557.get(0);
        mod_545.put(1, t);
    endrule
    rule rule_728;
        ChannelMessage t;
        t <- mod_539.get(0);
        mod_572.put(0, t);
    endrule
    rule rule_729;
        ChannelMessage t;
        t <- mod_541.get(1);
        mod_542.put(0, t);
    endrule
    rule rule_730;
        ChannelMessage t;
        t <- mod_555.get(0);
        mod_553.put(0, t);
    endrule
    rule rule_731;
        ChannelMessage t;
        t <- mod_567.get(0);
        mod_568.put(0, t);
    endrule
    rule rule_732;
        ChannelMessage t;
        t <- mod_535.get(0);
        mod_536.put(0, t);
    endrule
    rule rule_733;
        ChannelMessage t;
        t <- mod_549.get(0);
        mod_551.put(0, t);
    endrule
    rule rule_734;
        ChannelMessage t;
        t <- mod_552.get(0);
        mod_552.put(1, t);
    endrule
    rule rule_735;
        ChannelMessage t;
        t <- mod_553.get(1);
        mod_546.put(1, t);
    endrule
    rule rule_736;
        ChannelMessage t;
        t <- mod_562.get(0);
        mod_561.put(1, t);
    endrule
    rule rule_737;
        ChannelMessage t;
        t <- mod_561.get(1);
        mod_560.put(1, t);
    endrule
    rule rule_738;
        ChannelMessage t;
        t <- mod_563.get(0);
        mod_561.put(0, t);
    endrule
    rule rule_739;
        ChannelMessage t;
        t <- mod_548.get(0);
        mod_552.put(0, t);
    endrule
    rule rule_740;
        ChannelMessage t;
        t <- mod_545.get(1);
        mod_546.put(0, t);
    endrule
    rule rule_741;
        ChannelMessage t;
        t <- mod_567.get(1);
        mod_542.put(1, t);
    endrule
    rule rule_742;
        ChannelMessage t;
        t <- mod_538.get(3);
        mod_539.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_534.put(0, t);
        end
        if (i == 1) begin
            mod_550.put(0, t);
        end
        if (i == 2) begin
            mod_556.put(0, t);
        end
        if (i == 3) begin
            mod_564.put(0, t);
        end
        if (i == 4) begin
            mod_570.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_538.get(0);
        end
        if (i == 2) begin
            t <- mod_538.get(1);
        end
        if (i == 1) begin
            t <- mod_538.get(2);
        end
        if (i == 3) begin
            t <- mod_550.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6048 (Operation_IFC);
    Operation_IFC mod_575_inner <- mkReshape(2, 64);
    Operation_IFC mod_575 <- mkDebugOperation(mod_575_inner, "mod_575");
    Operation_IFC mod_576_inner <- mkFlatten(1);
    Operation_IFC mod_576 <- mkDebugOperation(mod_576_inner, "mod_576");
    Operation_IFC mod_577_inner <- mkFlatten(2);
    Operation_IFC mod_577 <- mkDebugOperation(mod_577_inner, "mod_577");
    Operation_IFC mod_578_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_578 <- mkDebugOperation(mod_578_inner, "mod_578");
    Broadcast_IFC#(4) mod_579_inner <- mkBroadcast(4);
    Operation_IFC mod_579 <- mkDebugOperation(mod_579_inner.op, "mod_579");
    PMU_IFC mod_580_bufferize <- mkPMU(2);
    Operation_IFC mod_580_inner = mod_580_bufferize.operation;
    Operation_IFC mod_580 <- mkDebugOperation(mod_580_inner, "mod_580");
    Broadcast_IFC#(2) mod_581_inner <- mkBroadcast(2);
    Operation_IFC mod_581 <- mkDebugOperation(mod_581_inner.op, "mod_581");
    PMU_IFC mod_582_bufferize <- mkPMU(1);
    Operation_IFC mod_582_inner = mod_582_bufferize.operation;
    Operation_IFC mod_582 <- mkDebugOperation(mod_582_inner, "mod_582");
    Operation_IFC mod_583_inner <- mkBinaryMap(1142, matmul_t_tile);
    Operation_IFC mod_583 <- mkDebugOperation(mod_583_inner, "mod_583");
    Operation_IFC mod_584_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_584 <- mkDebugOperation(mod_584_inner, "mod_584");
    Operation_IFC mod_585_inner <- mkBinaryMap(1910, mul_tile);
    Operation_IFC mod_585 <- mkDebugOperation(mod_585_inner, "mod_585");
    PMU_IFC mod_586_bufferize <- mkPMU(1);
    Operation_IFC mod_586_inner = mod_586_bufferize.operation;
    Operation_IFC mod_586 <- mkDebugOperation(mod_586_inner, "mod_586");
    Operation_IFC mod_587_inner <- mkBinaryMap(2535, matmul_t_tile);
    Operation_IFC mod_587 <- mkDebugOperation(mod_587_inner, "mod_587");
    Operation_IFC mod_588_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_588 <- mkDebugOperation(mod_588_inner, "mod_588");
    Operation_IFC mod_589_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_589 <- mkDebugOperation(mod_589_inner, "mod_589");
    Operation_IFC mod_590_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_590 <- mkDebugOperation(mod_590_inner, "mod_590");
    Operation_IFC mod_591_inner <- mkBinaryMap(2809, mul_tile);
    Operation_IFC mod_591 <- mkDebugOperation(mod_591_inner, "mod_591");
    PMU_IFC mod_592_bufferize <- mkPMU(1);
    Operation_IFC mod_592_inner = mod_592_bufferize.operation;
    Operation_IFC mod_592 <- mkDebugOperation(mod_592_inner, "mod_592");
    PMU_IFC mod_593_bufferize <- mkPMU(2);
    Operation_IFC mod_593_inner = mod_593_bufferize.operation;
    Operation_IFC mod_593 <- mkDebugOperation(mod_593_inner, "mod_593");
    PMU_IFC mod_594_bufferize <- mkPMU(2);
    Operation_IFC mod_594_inner = mod_594_bufferize.operation;
    Operation_IFC mod_594 <- mkDebugOperation(mod_594_inner, "mod_594");
    Operation_IFC mod_595_inner <- mkRepeatStatic(8);
    Operation_IFC mod_595 <- mkDebugOperation(mod_595_inner, "mod_595");
    Operation_IFC mod_596_inner <- mkFlatten(1);
    Operation_IFC mod_596 <- mkDebugOperation(mod_596_inner, "mod_596");
    Operation_IFC mod_597_inner <- mkFlatten(0);
    Operation_IFC mod_597 <- mkDebugOperation(mod_597_inner, "mod_597");
    Operation_IFC mod_598_inner <- mkRepeatStatic(3);
    Operation_IFC mod_598 <- mkDebugOperation(mod_598_inner, "mod_598");
    Operation_IFC mod_599_inner <- mkUnaryMap(1782, silu_tile);
    Operation_IFC mod_599 <- mkDebugOperation(mod_599_inner, "mod_599");
    Operation_IFC mod_600_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_600 <- mkDebugOperation(mod_600_inner, "mod_600");
    Operation_IFC mod_601_inner <- mkBinaryMap(1654, matmul_t_tile);
    Operation_IFC mod_601 <- mkDebugOperation(mod_601_inner, "mod_601");
    PMU_IFC mod_602_bufferize <- mkPMU(2);
    Operation_IFC mod_602_inner = mod_602_bufferize.operation;
    Operation_IFC mod_602 <- mkDebugOperation(mod_602_inner, "mod_602");
    Operation_IFC mod_603_inner <- mkRepeatStatic(8);
    Operation_IFC mod_603 <- mkDebugOperation(mod_603_inner, "mod_603");
    Operation_IFC mod_604_inner <- mkFlatten(1);
    Operation_IFC mod_604 <- mkDebugOperation(mod_604_inner, "mod_604");
    Operation_IFC mod_605_inner <- mkFlatten(0);
    Operation_IFC mod_605 <- mkDebugOperation(mod_605_inner, "mod_605");
    PMU_IFC mod_606_bufferize <- mkPMU(1);
    Operation_IFC mod_606_inner = mod_606_bufferize.operation;
    Operation_IFC mod_606 <- mkDebugOperation(mod_606_inner, "mod_606");
    Operation_IFC mod_607_inner <- mkRepeatStatic(16);
    Operation_IFC mod_607 <- mkDebugOperation(mod_607_inner, "mod_607");
    PMU_IFC mod_608_bufferize <- mkPMU(2);
    Operation_IFC mod_608_inner = mod_608_bufferize.operation;
    Operation_IFC mod_608 <- mkDebugOperation(mod_608_inner, "mod_608");
    Operation_IFC mod_609_inner <- mkRepeatStatic(8);
    Operation_IFC mod_609 <- mkDebugOperation(mod_609_inner, "mod_609");
    Operation_IFC mod_610_inner <- mkFlatten(1);
    Operation_IFC mod_610 <- mkDebugOperation(mod_610_inner, "mod_610");
    Operation_IFC mod_611_inner <- mkFlatten(0);
    Operation_IFC mod_611 <- mkDebugOperation(mod_611_inner, "mod_611");
    Operation_IFC mod_612_inner <- mkRepeatStatic(16);
    Operation_IFC mod_612 <- mkDebugOperation(mod_612_inner, "mod_612");
    Operation_IFC mod_613_inner <- mkRepeatStatic(2);
    Operation_IFC mod_613 <- mkDebugOperation(mod_613_inner, "mod_613");
    PMU_IFC mod_614_bufferize <- mkPMU(2);
    Operation_IFC mod_614_inner = mod_614_bufferize.operation;
    Operation_IFC mod_614 <- mkDebugOperation(mod_614_inner, "mod_614");
    rule rule_743;
        ChannelMessage t;
        t <- mod_592.get(1);
        mod_590.put(1, t);
    endrule
    rule rule_744;
        ChannelMessage t;
        t <- mod_602.get(0);
        mod_603.put(0, t);
    endrule
    rule rule_745;
        ChannelMessage t;
        t <- mod_605.get(0);
        mod_604.put(0, t);
    endrule
    rule rule_746;
        ChannelMessage t;
        t <- mod_612.get(0);
        mod_582.put(1, t);
    endrule
    rule rule_747;
        ChannelMessage t;
        t <- mod_584.get(0);
        mod_585.put(0, t);
    endrule
    rule rule_748;
        ChannelMessage t;
        t <- mod_578.get(1);
        mod_579.put(0, t);
    endrule
    rule rule_749;
        ChannelMessage t;
        t <- mod_596.get(0);
        mod_594.put(0, t);
    endrule
    rule rule_750;
        ChannelMessage t;
        t <- mod_608.get(1);
        mod_583.put(1, t);
    endrule
    rule rule_751;
        ChannelMessage t;
        t <- mod_609.get(0);
        mod_608.put(1, t);
    endrule
    rule rule_752;
        ChannelMessage t;
        t <- mod_590.get(0);
        mod_592.put(0, t);
    endrule
    rule rule_753;
        ChannelMessage t;
        t <- mod_610.get(0);
        mod_608.put(0, t);
    endrule
    rule rule_754;
        ChannelMessage t;
        t <- mod_580.get(0);
        mod_613.put(0, t);
    endrule
    rule rule_755;
        ChannelMessage t;
        t <- mod_590.get(1);
        mod_591.put(1, t);
    endrule
    rule rule_756;
        ChannelMessage t;
        t <- mod_597.get(0);
        mod_596.put(0, t);
    endrule
    rule rule_757;
        ChannelMessage t;
        t <- mod_581.get(1);
        mod_582.put(0, t);
    endrule
    rule rule_758;
        ChannelMessage t;
        t <- mod_588.get(0);
        mod_589.put(0, t);
    endrule
    rule rule_759;
        ChannelMessage t;
        t <- mod_580.get(1);
        mod_581.put(0, t);
    endrule
    rule rule_760;
        ChannelMessage t;
        t <- mod_575.get(0);
        mod_576.put(0, t);
    endrule
    rule rule_761;
        ChannelMessage t;
        t <- mod_586.get(0);
        mod_598.put(0, t);
    endrule
    rule rule_762;
        ChannelMessage t;
        t <- mod_585.get(0);
        mod_586.put(0, t);
    endrule
    rule rule_763;
        ChannelMessage t;
        t <- mod_606.get(1);
        mod_601.put(0, t);
    endrule
    rule rule_764;
        ChannelMessage t;
        t <- mod_586.get(1);
        mod_587.put(0, t);
    endrule
    rule rule_765;
        ChannelMessage t;
        t <- mod_595.get(0);
        mod_594.put(1, t);
    endrule
    rule rule_766;
        ChannelMessage t;
        t <- mod_601.get(0);
        mod_600.put(0, t);
    endrule
    rule rule_767;
        ChannelMessage t;
        t <- mod_611.get(0);
        mod_610.put(0, t);
    endrule
    rule rule_768;
        ChannelMessage t;
        t <- mod_587.get(0);
        mod_588.put(0, t);
    endrule
    rule rule_769;
        ChannelMessage t;
        t <- mod_578.get(0);
        mod_614.put(0, t);
    endrule
    rule rule_770;
        ChannelMessage t;
        t <- mod_589.get(1);
        mod_590.put(0, t);
    endrule
    rule rule_771;
        ChannelMessage t;
        t <- mod_599.get(0);
        mod_585.put(1, t);
    endrule
    rule rule_772;
        ChannelMessage t;
        t <- mod_579.get(3);
        mod_580.put(0, t);
    endrule
    rule rule_773;
        ChannelMessage t;
        t <- mod_608.get(0);
        mod_609.put(0, t);
    endrule
    rule rule_774;
        ChannelMessage t;
        t <- mod_602.get(1);
        mod_601.put(1, t);
    endrule
    rule rule_775;
        ChannelMessage t;
        t <- mod_593.get(1);
        mod_589.put(1, t);
    endrule
    rule rule_776;
        ChannelMessage t;
        t <- mod_603.get(0);
        mod_602.put(1, t);
    endrule
    rule rule_777;
        ChannelMessage t;
        t <- mod_604.get(0);
        mod_602.put(0, t);
    endrule
    rule rule_778;
        ChannelMessage t;
        t <- mod_577.get(0);
        mod_578.put(0, t);
    endrule
    rule rule_779;
        ChannelMessage t;
        t <- mod_594.get(0);
        mod_595.put(0, t);
    endrule
    rule rule_780;
        ChannelMessage t;
        t <- mod_607.get(0);
        mod_606.put(1, t);
    endrule
    rule rule_781;
        ChannelMessage t;
        t <- mod_589.get(0);
        mod_593.put(0, t);
    endrule
    rule rule_782;
        ChannelMessage t;
        t <- mod_592.get(0);
        mod_592.put(1, t);
    endrule
    rule rule_783;
        ChannelMessage t;
        t <- mod_614.get(0);
        mod_614.put(1, t);
    endrule
    rule rule_784;
        ChannelMessage t;
        t <- mod_593.get(0);
        mod_593.put(1, t);
    endrule
    rule rule_785;
        ChannelMessage t;
        t <- mod_613.get(0);
        mod_580.put(1, t);
    endrule
    rule rule_786;
        ChannelMessage t;
        t <- mod_582.get(0);
        mod_612.put(0, t);
    endrule
    rule rule_787;
        ChannelMessage t;
        t <- mod_614.get(1);
        mod_578.put(1, t);
    endrule
    rule rule_788;
        ChannelMessage t;
        t <- mod_582.get(1);
        mod_583.put(0, t);
    endrule
    rule rule_789;
        ChannelMessage t;
        t <- mod_606.get(0);
        mod_607.put(0, t);
    endrule
    rule rule_790;
        ChannelMessage t;
        t <- mod_576.get(0);
        mod_577.put(0, t);
    endrule
    rule rule_791;
        ChannelMessage t;
        t <- mod_583.get(0);
        mod_584.put(0, t);
    endrule
    rule rule_792;
        ChannelMessage t;
        t <- mod_594.get(1);
        mod_587.put(1, t);
    endrule
    rule rule_793;
        ChannelMessage t;
        t <- mod_600.get(0);
        mod_599.put(0, t);
    endrule
    rule rule_794;
        ChannelMessage t;
        t <- mod_581.get(0);
        mod_606.put(0, t);
    endrule
    rule rule_795;
        ChannelMessage t;
        t <- mod_598.get(0);
        mod_586.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_575.put(0, t);
        end
        if (i == 1) begin
            mod_591.put(0, t);
        end
        if (i == 2) begin
            mod_597.put(0, t);
        end
        if (i == 3) begin
            mod_605.put(0, t);
        end
        if (i == 4) begin
            mod_611.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_579.get(0);
        end
        if (i == 2) begin
            t <- mod_579.get(1);
        end
        if (i == 3) begin
            t <- mod_579.get(2);
        end
        if (i == 1) begin
            t <- mod_591.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6049 (Operation_IFC);
    Operation_IFC mod_616_inner <- mkReshape(2, 64);
    Operation_IFC mod_616 <- mkDebugOperation(mod_616_inner, "mod_616");
    Operation_IFC mod_617_inner <- mkFlatten(1);
    Operation_IFC mod_617 <- mkDebugOperation(mod_617_inner, "mod_617");
    Operation_IFC mod_618_inner <- mkFlatten(2);
    Operation_IFC mod_618 <- mkDebugOperation(mod_618_inner, "mod_618");
    Operation_IFC mod_619_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_619 <- mkDebugOperation(mod_619_inner, "mod_619");
    Broadcast_IFC#(4) mod_620_inner <- mkBroadcast(4);
    Operation_IFC mod_620 <- mkDebugOperation(mod_620_inner.op, "mod_620");
    PMU_IFC mod_621_bufferize <- mkPMU(2);
    Operation_IFC mod_621_inner = mod_621_bufferize.operation;
    Operation_IFC mod_621 <- mkDebugOperation(mod_621_inner, "mod_621");
    Broadcast_IFC#(2) mod_622_inner <- mkBroadcast(2);
    Operation_IFC mod_622 <- mkDebugOperation(mod_622_inner.op, "mod_622");
    PMU_IFC mod_623_bufferize <- mkPMU(1);
    Operation_IFC mod_623_inner = mod_623_bufferize.operation;
    Operation_IFC mod_623 <- mkDebugOperation(mod_623_inner, "mod_623");
    Operation_IFC mod_624_inner <- mkBinaryMap(1141, matmul_t_tile);
    Operation_IFC mod_624 <- mkDebugOperation(mod_624_inner, "mod_624");
    Operation_IFC mod_625_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_625 <- mkDebugOperation(mod_625_inner, "mod_625");
    Operation_IFC mod_626_inner <- mkBinaryMap(1909, mul_tile);
    Operation_IFC mod_626 <- mkDebugOperation(mod_626_inner, "mod_626");
    PMU_IFC mod_627_bufferize <- mkPMU(1);
    Operation_IFC mod_627_inner = mod_627_bufferize.operation;
    Operation_IFC mod_627 <- mkDebugOperation(mod_627_inner, "mod_627");
    Operation_IFC mod_628_inner <- mkBinaryMap(2533, matmul_t_tile);
    Operation_IFC mod_628 <- mkDebugOperation(mod_628_inner, "mod_628");
    Operation_IFC mod_629_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_629 <- mkDebugOperation(mod_629_inner, "mod_629");
    Operation_IFC mod_630_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_630 <- mkDebugOperation(mod_630_inner, "mod_630");
    Operation_IFC mod_631_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_631 <- mkDebugOperation(mod_631_inner, "mod_631");
    Operation_IFC mod_632_inner <- mkBinaryMap(2808, mul_tile);
    Operation_IFC mod_632 <- mkDebugOperation(mod_632_inner, "mod_632");
    PMU_IFC mod_633_bufferize <- mkPMU(1);
    Operation_IFC mod_633_inner = mod_633_bufferize.operation;
    Operation_IFC mod_633 <- mkDebugOperation(mod_633_inner, "mod_633");
    PMU_IFC mod_634_bufferize <- mkPMU(2);
    Operation_IFC mod_634_inner = mod_634_bufferize.operation;
    Operation_IFC mod_634 <- mkDebugOperation(mod_634_inner, "mod_634");
    PMU_IFC mod_635_bufferize <- mkPMU(2);
    Operation_IFC mod_635_inner = mod_635_bufferize.operation;
    Operation_IFC mod_635 <- mkDebugOperation(mod_635_inner, "mod_635");
    Operation_IFC mod_636_inner <- mkRepeatStatic(8);
    Operation_IFC mod_636 <- mkDebugOperation(mod_636_inner, "mod_636");
    Operation_IFC mod_637_inner <- mkFlatten(1);
    Operation_IFC mod_637 <- mkDebugOperation(mod_637_inner, "mod_637");
    Operation_IFC mod_638_inner <- mkFlatten(0);
    Operation_IFC mod_638 <- mkDebugOperation(mod_638_inner, "mod_638");
    Operation_IFC mod_639_inner <- mkRepeatStatic(3);
    Operation_IFC mod_639 <- mkDebugOperation(mod_639_inner, "mod_639");
    Operation_IFC mod_640_inner <- mkUnaryMap(1781, silu_tile);
    Operation_IFC mod_640 <- mkDebugOperation(mod_640_inner, "mod_640");
    Operation_IFC mod_641_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_641 <- mkDebugOperation(mod_641_inner, "mod_641");
    Operation_IFC mod_642_inner <- mkBinaryMap(1653, matmul_t_tile);
    Operation_IFC mod_642 <- mkDebugOperation(mod_642_inner, "mod_642");
    PMU_IFC mod_643_bufferize <- mkPMU(2);
    Operation_IFC mod_643_inner = mod_643_bufferize.operation;
    Operation_IFC mod_643 <- mkDebugOperation(mod_643_inner, "mod_643");
    Operation_IFC mod_644_inner <- mkRepeatStatic(8);
    Operation_IFC mod_644 <- mkDebugOperation(mod_644_inner, "mod_644");
    Operation_IFC mod_645_inner <- mkFlatten(1);
    Operation_IFC mod_645 <- mkDebugOperation(mod_645_inner, "mod_645");
    Operation_IFC mod_646_inner <- mkFlatten(0);
    Operation_IFC mod_646 <- mkDebugOperation(mod_646_inner, "mod_646");
    PMU_IFC mod_647_bufferize <- mkPMU(1);
    Operation_IFC mod_647_inner = mod_647_bufferize.operation;
    Operation_IFC mod_647 <- mkDebugOperation(mod_647_inner, "mod_647");
    Operation_IFC mod_648_inner <- mkRepeatStatic(16);
    Operation_IFC mod_648 <- mkDebugOperation(mod_648_inner, "mod_648");
    PMU_IFC mod_649_bufferize <- mkPMU(2);
    Operation_IFC mod_649_inner = mod_649_bufferize.operation;
    Operation_IFC mod_649 <- mkDebugOperation(mod_649_inner, "mod_649");
    Operation_IFC mod_650_inner <- mkRepeatStatic(8);
    Operation_IFC mod_650 <- mkDebugOperation(mod_650_inner, "mod_650");
    Operation_IFC mod_651_inner <- mkFlatten(1);
    Operation_IFC mod_651 <- mkDebugOperation(mod_651_inner, "mod_651");
    Operation_IFC mod_652_inner <- mkFlatten(0);
    Operation_IFC mod_652 <- mkDebugOperation(mod_652_inner, "mod_652");
    Operation_IFC mod_653_inner <- mkRepeatStatic(16);
    Operation_IFC mod_653 <- mkDebugOperation(mod_653_inner, "mod_653");
    Operation_IFC mod_654_inner <- mkRepeatStatic(2);
    Operation_IFC mod_654 <- mkDebugOperation(mod_654_inner, "mod_654");
    PMU_IFC mod_655_bufferize <- mkPMU(2);
    Operation_IFC mod_655_inner = mod_655_bufferize.operation;
    Operation_IFC mod_655 <- mkDebugOperation(mod_655_inner, "mod_655");
    rule rule_796;
        ChannelMessage t;
        t <- mod_626.get(0);
        mod_627.put(0, t);
    endrule
    rule rule_797;
        ChannelMessage t;
        t <- mod_623.get(1);
        mod_624.put(0, t);
    endrule
    rule rule_798;
        ChannelMessage t;
        t <- mod_637.get(0);
        mod_635.put(0, t);
    endrule
    rule rule_799;
        ChannelMessage t;
        t <- mod_645.get(0);
        mod_643.put(0, t);
    endrule
    rule rule_800;
        ChannelMessage t;
        t <- mod_630.get(0);
        mod_634.put(0, t);
    endrule
    rule rule_801;
        ChannelMessage t;
        t <- mod_654.get(0);
        mod_621.put(1, t);
    endrule
    rule rule_802;
        ChannelMessage t;
        t <- mod_635.get(1);
        mod_628.put(1, t);
    endrule
    rule rule_803;
        ChannelMessage t;
        t <- mod_650.get(0);
        mod_649.put(1, t);
    endrule
    rule rule_804;
        ChannelMessage t;
        t <- mod_646.get(0);
        mod_645.put(0, t);
    endrule
    rule rule_805;
        ChannelMessage t;
        t <- mod_655.get(1);
        mod_619.put(1, t);
    endrule
    rule rule_806;
        ChannelMessage t;
        t <- mod_643.get(0);
        mod_644.put(0, t);
    endrule
    rule rule_807;
        ChannelMessage t;
        t <- mod_639.get(0);
        mod_627.put(1, t);
    endrule
    rule rule_808;
        ChannelMessage t;
        t <- mod_647.get(1);
        mod_642.put(0, t);
    endrule
    rule rule_809;
        ChannelMessage t;
        t <- mod_616.get(0);
        mod_617.put(0, t);
    endrule
    rule rule_810;
        ChannelMessage t;
        t <- mod_634.get(0);
        mod_634.put(1, t);
    endrule
    rule rule_811;
        ChannelMessage t;
        t <- mod_617.get(0);
        mod_618.put(0, t);
    endrule
    rule rule_812;
        ChannelMessage t;
        t <- mod_653.get(0);
        mod_623.put(1, t);
    endrule
    rule rule_813;
        ChannelMessage t;
        t <- mod_623.get(0);
        mod_653.put(0, t);
    endrule
    rule rule_814;
        ChannelMessage t;
        t <- mod_630.get(1);
        mod_631.put(0, t);
    endrule
    rule rule_815;
        ChannelMessage t;
        t <- mod_643.get(1);
        mod_642.put(1, t);
    endrule
    rule rule_816;
        ChannelMessage t;
        t <- mod_635.get(0);
        mod_636.put(0, t);
    endrule
    rule rule_817;
        ChannelMessage t;
        t <- mod_619.get(0);
        mod_655.put(0, t);
    endrule
    rule rule_818;
        ChannelMessage t;
        t <- mod_649.get(1);
        mod_624.put(1, t);
    endrule
    rule rule_819;
        ChannelMessage t;
        t <- mod_621.get(1);
        mod_622.put(0, t);
    endrule
    rule rule_820;
        ChannelMessage t;
        t <- mod_631.get(1);
        mod_632.put(1, t);
    endrule
    rule rule_821;
        ChannelMessage t;
        t <- mod_641.get(0);
        mod_640.put(0, t);
    endrule
    rule rule_822;
        ChannelMessage t;
        t <- mod_619.get(1);
        mod_620.put(0, t);
    endrule
    rule rule_823;
        ChannelMessage t;
        t <- mod_621.get(0);
        mod_654.put(0, t);
    endrule
    rule rule_824;
        ChannelMessage t;
        t <- mod_627.get(0);
        mod_639.put(0, t);
    endrule
    rule rule_825;
        ChannelMessage t;
        t <- mod_624.get(0);
        mod_625.put(0, t);
    endrule
    rule rule_826;
        ChannelMessage t;
        t <- mod_634.get(1);
        mod_630.put(1, t);
    endrule
    rule rule_827;
        ChannelMessage t;
        t <- mod_622.get(0);
        mod_647.put(0, t);
    endrule
    rule rule_828;
        ChannelMessage t;
        t <- mod_644.get(0);
        mod_643.put(1, t);
    endrule
    rule rule_829;
        ChannelMessage t;
        t <- mod_652.get(0);
        mod_651.put(0, t);
    endrule
    rule rule_830;
        ChannelMessage t;
        t <- mod_647.get(0);
        mod_648.put(0, t);
    endrule
    rule rule_831;
        ChannelMessage t;
        t <- mod_638.get(0);
        mod_637.put(0, t);
    endrule
    rule rule_832;
        ChannelMessage t;
        t <- mod_629.get(0);
        mod_630.put(0, t);
    endrule
    rule rule_833;
        ChannelMessage t;
        t <- mod_625.get(0);
        mod_626.put(0, t);
    endrule
    rule rule_834;
        ChannelMessage t;
        t <- mod_618.get(0);
        mod_619.put(0, t);
    endrule
    rule rule_835;
        ChannelMessage t;
        t <- mod_622.get(1);
        mod_623.put(0, t);
    endrule
    rule rule_836;
        ChannelMessage t;
        t <- mod_633.get(1);
        mod_631.put(1, t);
    endrule
    rule rule_837;
        ChannelMessage t;
        t <- mod_651.get(0);
        mod_649.put(0, t);
    endrule
    rule rule_838;
        ChannelMessage t;
        t <- mod_649.get(0);
        mod_650.put(0, t);
    endrule
    rule rule_839;
        ChannelMessage t;
        t <- mod_627.get(1);
        mod_628.put(0, t);
    endrule
    rule rule_840;
        ChannelMessage t;
        t <- mod_620.get(3);
        mod_621.put(0, t);
    endrule
    rule rule_841;
        ChannelMessage t;
        t <- mod_640.get(0);
        mod_626.put(1, t);
    endrule
    rule rule_842;
        ChannelMessage t;
        t <- mod_642.get(0);
        mod_641.put(0, t);
    endrule
    rule rule_843;
        ChannelMessage t;
        t <- mod_631.get(0);
        mod_633.put(0, t);
    endrule
    rule rule_844;
        ChannelMessage t;
        t <- mod_648.get(0);
        mod_647.put(1, t);
    endrule
    rule rule_845;
        ChannelMessage t;
        t <- mod_628.get(0);
        mod_629.put(0, t);
    endrule
    rule rule_846;
        ChannelMessage t;
        t <- mod_655.get(0);
        mod_655.put(1, t);
    endrule
    rule rule_847;
        ChannelMessage t;
        t <- mod_636.get(0);
        mod_635.put(1, t);
    endrule
    rule rule_848;
        ChannelMessage t;
        t <- mod_633.get(0);
        mod_633.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_616.put(0, t);
        end
        if (i == 1) begin
            mod_632.put(0, t);
        end
        if (i == 2) begin
            mod_638.put(0, t);
        end
        if (i == 3) begin
            mod_646.put(0, t);
        end
        if (i == 4) begin
            mod_652.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_620.get(0);
        end
        if (i == 1) begin
            t <- mod_620.get(1);
        end
        if (i == 2) begin
            t <- mod_620.get(2);
        end
        if (i == 3) begin
            t <- mod_632.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6050 (Operation_IFC);
    Operation_IFC mod_657_inner <- mkReshape(2, 64);
    Operation_IFC mod_657 <- mkDebugOperation(mod_657_inner, "mod_657");
    Operation_IFC mod_658_inner <- mkFlatten(1);
    Operation_IFC mod_658 <- mkDebugOperation(mod_658_inner, "mod_658");
    Operation_IFC mod_659_inner <- mkFlatten(2);
    Operation_IFC mod_659 <- mkDebugOperation(mod_659_inner, "mod_659");
    Operation_IFC mod_660_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_660 <- mkDebugOperation(mod_660_inner, "mod_660");
    Broadcast_IFC#(4) mod_661_inner <- mkBroadcast(4);
    Operation_IFC mod_661 <- mkDebugOperation(mod_661_inner.op, "mod_661");
    PMU_IFC mod_662_bufferize <- mkPMU(2);
    Operation_IFC mod_662_inner = mod_662_bufferize.operation;
    Operation_IFC mod_662 <- mkDebugOperation(mod_662_inner, "mod_662");
    Broadcast_IFC#(2) mod_663_inner <- mkBroadcast(2);
    Operation_IFC mod_663 <- mkDebugOperation(mod_663_inner.op, "mod_663");
    PMU_IFC mod_664_bufferize <- mkPMU(1);
    Operation_IFC mod_664_inner = mod_664_bufferize.operation;
    Operation_IFC mod_664 <- mkDebugOperation(mod_664_inner, "mod_664");
    Operation_IFC mod_665_inner <- mkBinaryMap(1140, matmul_t_tile);
    Operation_IFC mod_665 <- mkDebugOperation(mod_665_inner, "mod_665");
    Operation_IFC mod_666_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_666 <- mkDebugOperation(mod_666_inner, "mod_666");
    Operation_IFC mod_667_inner <- mkBinaryMap(1908, mul_tile);
    Operation_IFC mod_667 <- mkDebugOperation(mod_667_inner, "mod_667");
    PMU_IFC mod_668_bufferize <- mkPMU(1);
    Operation_IFC mod_668_inner = mod_668_bufferize.operation;
    Operation_IFC mod_668 <- mkDebugOperation(mod_668_inner, "mod_668");
    Operation_IFC mod_669_inner <- mkBinaryMap(2531, matmul_t_tile);
    Operation_IFC mod_669 <- mkDebugOperation(mod_669_inner, "mod_669");
    Operation_IFC mod_670_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_670 <- mkDebugOperation(mod_670_inner, "mod_670");
    Operation_IFC mod_671_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_671 <- mkDebugOperation(mod_671_inner, "mod_671");
    Operation_IFC mod_672_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_672 <- mkDebugOperation(mod_672_inner, "mod_672");
    Operation_IFC mod_673_inner <- mkBinaryMap(2807, mul_tile);
    Operation_IFC mod_673 <- mkDebugOperation(mod_673_inner, "mod_673");
    PMU_IFC mod_674_bufferize <- mkPMU(1);
    Operation_IFC mod_674_inner = mod_674_bufferize.operation;
    Operation_IFC mod_674 <- mkDebugOperation(mod_674_inner, "mod_674");
    PMU_IFC mod_675_bufferize <- mkPMU(2);
    Operation_IFC mod_675_inner = mod_675_bufferize.operation;
    Operation_IFC mod_675 <- mkDebugOperation(mod_675_inner, "mod_675");
    PMU_IFC mod_676_bufferize <- mkPMU(2);
    Operation_IFC mod_676_inner = mod_676_bufferize.operation;
    Operation_IFC mod_676 <- mkDebugOperation(mod_676_inner, "mod_676");
    Operation_IFC mod_677_inner <- mkRepeatStatic(8);
    Operation_IFC mod_677 <- mkDebugOperation(mod_677_inner, "mod_677");
    Operation_IFC mod_678_inner <- mkFlatten(1);
    Operation_IFC mod_678 <- mkDebugOperation(mod_678_inner, "mod_678");
    Operation_IFC mod_679_inner <- mkFlatten(0);
    Operation_IFC mod_679 <- mkDebugOperation(mod_679_inner, "mod_679");
    Operation_IFC mod_680_inner <- mkRepeatStatic(3);
    Operation_IFC mod_680 <- mkDebugOperation(mod_680_inner, "mod_680");
    Operation_IFC mod_681_inner <- mkUnaryMap(1780, silu_tile);
    Operation_IFC mod_681 <- mkDebugOperation(mod_681_inner, "mod_681");
    Operation_IFC mod_682_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_682 <- mkDebugOperation(mod_682_inner, "mod_682");
    Operation_IFC mod_683_inner <- mkBinaryMap(1652, matmul_t_tile);
    Operation_IFC mod_683 <- mkDebugOperation(mod_683_inner, "mod_683");
    PMU_IFC mod_684_bufferize <- mkPMU(2);
    Operation_IFC mod_684_inner = mod_684_bufferize.operation;
    Operation_IFC mod_684 <- mkDebugOperation(mod_684_inner, "mod_684");
    Operation_IFC mod_685_inner <- mkRepeatStatic(8);
    Operation_IFC mod_685 <- mkDebugOperation(mod_685_inner, "mod_685");
    Operation_IFC mod_686_inner <- mkFlatten(1);
    Operation_IFC mod_686 <- mkDebugOperation(mod_686_inner, "mod_686");
    Operation_IFC mod_687_inner <- mkFlatten(0);
    Operation_IFC mod_687 <- mkDebugOperation(mod_687_inner, "mod_687");
    PMU_IFC mod_688_bufferize <- mkPMU(1);
    Operation_IFC mod_688_inner = mod_688_bufferize.operation;
    Operation_IFC mod_688 <- mkDebugOperation(mod_688_inner, "mod_688");
    Operation_IFC mod_689_inner <- mkRepeatStatic(16);
    Operation_IFC mod_689 <- mkDebugOperation(mod_689_inner, "mod_689");
    PMU_IFC mod_690_bufferize <- mkPMU(2);
    Operation_IFC mod_690_inner = mod_690_bufferize.operation;
    Operation_IFC mod_690 <- mkDebugOperation(mod_690_inner, "mod_690");
    Operation_IFC mod_691_inner <- mkRepeatStatic(8);
    Operation_IFC mod_691 <- mkDebugOperation(mod_691_inner, "mod_691");
    Operation_IFC mod_692_inner <- mkFlatten(1);
    Operation_IFC mod_692 <- mkDebugOperation(mod_692_inner, "mod_692");
    Operation_IFC mod_693_inner <- mkFlatten(0);
    Operation_IFC mod_693 <- mkDebugOperation(mod_693_inner, "mod_693");
    Operation_IFC mod_694_inner <- mkRepeatStatic(16);
    Operation_IFC mod_694 <- mkDebugOperation(mod_694_inner, "mod_694");
    Operation_IFC mod_695_inner <- mkRepeatStatic(2);
    Operation_IFC mod_695 <- mkDebugOperation(mod_695_inner, "mod_695");
    PMU_IFC mod_696_bufferize <- mkPMU(2);
    Operation_IFC mod_696_inner = mod_696_bufferize.operation;
    Operation_IFC mod_696 <- mkDebugOperation(mod_696_inner, "mod_696");
    rule rule_849;
        ChannelMessage t;
        t <- mod_663.get(0);
        mod_688.put(0, t);
    endrule
    rule rule_850;
        ChannelMessage t;
        t <- mod_674.get(0);
        mod_674.put(1, t);
    endrule
    rule rule_851;
        ChannelMessage t;
        t <- mod_668.get(1);
        mod_669.put(0, t);
    endrule
    rule rule_852;
        ChannelMessage t;
        t <- mod_694.get(0);
        mod_664.put(1, t);
    endrule
    rule rule_853;
        ChannelMessage t;
        t <- mod_696.get(1);
        mod_660.put(1, t);
    endrule
    rule rule_854;
        ChannelMessage t;
        t <- mod_661.get(3);
        mod_662.put(0, t);
    endrule
    rule rule_855;
        ChannelMessage t;
        t <- mod_664.get(1);
        mod_665.put(0, t);
    endrule
    rule rule_856;
        ChannelMessage t;
        t <- mod_683.get(0);
        mod_682.put(0, t);
    endrule
    rule rule_857;
        ChannelMessage t;
        t <- mod_660.get(0);
        mod_696.put(0, t);
    endrule
    rule rule_858;
        ChannelMessage t;
        t <- mod_675.get(0);
        mod_675.put(1, t);
    endrule
    rule rule_859;
        ChannelMessage t;
        t <- mod_662.get(0);
        mod_695.put(0, t);
    endrule
    rule rule_860;
        ChannelMessage t;
        t <- mod_669.get(0);
        mod_670.put(0, t);
    endrule
    rule rule_861;
        ChannelMessage t;
        t <- mod_670.get(0);
        mod_671.put(0, t);
    endrule
    rule rule_862;
        ChannelMessage t;
        t <- mod_680.get(0);
        mod_668.put(1, t);
    endrule
    rule rule_863;
        ChannelMessage t;
        t <- mod_676.get(1);
        mod_669.put(1, t);
    endrule
    rule rule_864;
        ChannelMessage t;
        t <- mod_666.get(0);
        mod_667.put(0, t);
    endrule
    rule rule_865;
        ChannelMessage t;
        t <- mod_657.get(0);
        mod_658.put(0, t);
    endrule
    rule rule_866;
        ChannelMessage t;
        t <- mod_679.get(0);
        mod_678.put(0, t);
    endrule
    rule rule_867;
        ChannelMessage t;
        t <- mod_682.get(0);
        mod_681.put(0, t);
    endrule
    rule rule_868;
        ChannelMessage t;
        t <- mod_684.get(0);
        mod_685.put(0, t);
    endrule
    rule rule_869;
        ChannelMessage t;
        t <- mod_672.get(1);
        mod_673.put(1, t);
    endrule
    rule rule_870;
        ChannelMessage t;
        t <- mod_668.get(0);
        mod_680.put(0, t);
    endrule
    rule rule_871;
        ChannelMessage t;
        t <- mod_687.get(0);
        mod_686.put(0, t);
    endrule
    rule rule_872;
        ChannelMessage t;
        t <- mod_690.get(1);
        mod_665.put(1, t);
    endrule
    rule rule_873;
        ChannelMessage t;
        t <- mod_685.get(0);
        mod_684.put(1, t);
    endrule
    rule rule_874;
        ChannelMessage t;
        t <- mod_663.get(1);
        mod_664.put(0, t);
    endrule
    rule rule_875;
        ChannelMessage t;
        t <- mod_665.get(0);
        mod_666.put(0, t);
    endrule
    rule rule_876;
        ChannelMessage t;
        t <- mod_672.get(0);
        mod_674.put(0, t);
    endrule
    rule rule_877;
        ChannelMessage t;
        t <- mod_677.get(0);
        mod_676.put(1, t);
    endrule
    rule rule_878;
        ChannelMessage t;
        t <- mod_691.get(0);
        mod_690.put(1, t);
    endrule
    rule rule_879;
        ChannelMessage t;
        t <- mod_692.get(0);
        mod_690.put(0, t);
    endrule
    rule rule_880;
        ChannelMessage t;
        t <- mod_696.get(0);
        mod_696.put(1, t);
    endrule
    rule rule_881;
        ChannelMessage t;
        t <- mod_695.get(0);
        mod_662.put(1, t);
    endrule
    rule rule_882;
        ChannelMessage t;
        t <- mod_659.get(0);
        mod_660.put(0, t);
    endrule
    rule rule_883;
        ChannelMessage t;
        t <- mod_660.get(1);
        mod_661.put(0, t);
    endrule
    rule rule_884;
        ChannelMessage t;
        t <- mod_671.get(1);
        mod_672.put(0, t);
    endrule
    rule rule_885;
        ChannelMessage t;
        t <- mod_686.get(0);
        mod_684.put(0, t);
    endrule
    rule rule_886;
        ChannelMessage t;
        t <- mod_689.get(0);
        mod_688.put(1, t);
    endrule
    rule rule_887;
        ChannelMessage t;
        t <- mod_671.get(0);
        mod_675.put(0, t);
    endrule
    rule rule_888;
        ChannelMessage t;
        t <- mod_676.get(0);
        mod_677.put(0, t);
    endrule
    rule rule_889;
        ChannelMessage t;
        t <- mod_658.get(0);
        mod_659.put(0, t);
    endrule
    rule rule_890;
        ChannelMessage t;
        t <- mod_678.get(0);
        mod_676.put(0, t);
    endrule
    rule rule_891;
        ChannelMessage t;
        t <- mod_675.get(1);
        mod_671.put(1, t);
    endrule
    rule rule_892;
        ChannelMessage t;
        t <- mod_674.get(1);
        mod_672.put(1, t);
    endrule
    rule rule_893;
        ChannelMessage t;
        t <- mod_662.get(1);
        mod_663.put(0, t);
    endrule
    rule rule_894;
        ChannelMessage t;
        t <- mod_688.get(1);
        mod_683.put(0, t);
    endrule
    rule rule_895;
        ChannelMessage t;
        t <- mod_681.get(0);
        mod_667.put(1, t);
    endrule
    rule rule_896;
        ChannelMessage t;
        t <- mod_688.get(0);
        mod_689.put(0, t);
    endrule
    rule rule_897;
        ChannelMessage t;
        t <- mod_684.get(1);
        mod_683.put(1, t);
    endrule
    rule rule_898;
        ChannelMessage t;
        t <- mod_690.get(0);
        mod_691.put(0, t);
    endrule
    rule rule_899;
        ChannelMessage t;
        t <- mod_664.get(0);
        mod_694.put(0, t);
    endrule
    rule rule_900;
        ChannelMessage t;
        t <- mod_667.get(0);
        mod_668.put(0, t);
    endrule
    rule rule_901;
        ChannelMessage t;
        t <- mod_693.get(0);
        mod_692.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_657.put(0, t);
        end
        if (i == 1) begin
            mod_673.put(0, t);
        end
        if (i == 2) begin
            mod_679.put(0, t);
        end
        if (i == 3) begin
            mod_687.put(0, t);
        end
        if (i == 4) begin
            mod_693.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_661.get(0);
        end
        if (i == 0) begin
            t <- mod_661.get(1);
        end
        if (i == 2) begin
            t <- mod_661.get(2);
        end
        if (i == 3) begin
            t <- mod_673.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6051 (Operation_IFC);
    Operation_IFC mod_698_inner <- mkReshape(2, 64);
    Operation_IFC mod_698 <- mkDebugOperation(mod_698_inner, "mod_698");
    Operation_IFC mod_699_inner <- mkFlatten(1);
    Operation_IFC mod_699 <- mkDebugOperation(mod_699_inner, "mod_699");
    Operation_IFC mod_700_inner <- mkFlatten(2);
    Operation_IFC mod_700 <- mkDebugOperation(mod_700_inner, "mod_700");
    Operation_IFC mod_701_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_701 <- mkDebugOperation(mod_701_inner, "mod_701");
    Broadcast_IFC#(4) mod_702_inner <- mkBroadcast(4);
    Operation_IFC mod_702 <- mkDebugOperation(mod_702_inner.op, "mod_702");
    PMU_IFC mod_703_bufferize <- mkPMU(2);
    Operation_IFC mod_703_inner = mod_703_bufferize.operation;
    Operation_IFC mod_703 <- mkDebugOperation(mod_703_inner, "mod_703");
    Broadcast_IFC#(2) mod_704_inner <- mkBroadcast(2);
    Operation_IFC mod_704 <- mkDebugOperation(mod_704_inner.op, "mod_704");
    PMU_IFC mod_705_bufferize <- mkPMU(1);
    Operation_IFC mod_705_inner = mod_705_bufferize.operation;
    Operation_IFC mod_705 <- mkDebugOperation(mod_705_inner, "mod_705");
    Operation_IFC mod_706_inner <- mkBinaryMap(1139, matmul_t_tile);
    Operation_IFC mod_706 <- mkDebugOperation(mod_706_inner, "mod_706");
    Operation_IFC mod_707_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_707 <- mkDebugOperation(mod_707_inner, "mod_707");
    Operation_IFC mod_708_inner <- mkBinaryMap(1907, mul_tile);
    Operation_IFC mod_708 <- mkDebugOperation(mod_708_inner, "mod_708");
    PMU_IFC mod_709_bufferize <- mkPMU(1);
    Operation_IFC mod_709_inner = mod_709_bufferize.operation;
    Operation_IFC mod_709 <- mkDebugOperation(mod_709_inner, "mod_709");
    Operation_IFC mod_710_inner <- mkBinaryMap(2529, matmul_t_tile);
    Operation_IFC mod_710 <- mkDebugOperation(mod_710_inner, "mod_710");
    Operation_IFC mod_711_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_711 <- mkDebugOperation(mod_711_inner, "mod_711");
    Operation_IFC mod_712_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_712 <- mkDebugOperation(mod_712_inner, "mod_712");
    Operation_IFC mod_713_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_713 <- mkDebugOperation(mod_713_inner, "mod_713");
    Operation_IFC mod_714_inner <- mkBinaryMap(2806, mul_tile);
    Operation_IFC mod_714 <- mkDebugOperation(mod_714_inner, "mod_714");
    PMU_IFC mod_715_bufferize <- mkPMU(1);
    Operation_IFC mod_715_inner = mod_715_bufferize.operation;
    Operation_IFC mod_715 <- mkDebugOperation(mod_715_inner, "mod_715");
    PMU_IFC mod_716_bufferize <- mkPMU(2);
    Operation_IFC mod_716_inner = mod_716_bufferize.operation;
    Operation_IFC mod_716 <- mkDebugOperation(mod_716_inner, "mod_716");
    PMU_IFC mod_717_bufferize <- mkPMU(2);
    Operation_IFC mod_717_inner = mod_717_bufferize.operation;
    Operation_IFC mod_717 <- mkDebugOperation(mod_717_inner, "mod_717");
    Operation_IFC mod_718_inner <- mkRepeatStatic(8);
    Operation_IFC mod_718 <- mkDebugOperation(mod_718_inner, "mod_718");
    Operation_IFC mod_719_inner <- mkFlatten(1);
    Operation_IFC mod_719 <- mkDebugOperation(mod_719_inner, "mod_719");
    Operation_IFC mod_720_inner <- mkFlatten(0);
    Operation_IFC mod_720 <- mkDebugOperation(mod_720_inner, "mod_720");
    Operation_IFC mod_721_inner <- mkRepeatStatic(3);
    Operation_IFC mod_721 <- mkDebugOperation(mod_721_inner, "mod_721");
    Operation_IFC mod_722_inner <- mkUnaryMap(1779, silu_tile);
    Operation_IFC mod_722 <- mkDebugOperation(mod_722_inner, "mod_722");
    Operation_IFC mod_723_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_723 <- mkDebugOperation(mod_723_inner, "mod_723");
    Operation_IFC mod_724_inner <- mkBinaryMap(1651, matmul_t_tile);
    Operation_IFC mod_724 <- mkDebugOperation(mod_724_inner, "mod_724");
    PMU_IFC mod_725_bufferize <- mkPMU(2);
    Operation_IFC mod_725_inner = mod_725_bufferize.operation;
    Operation_IFC mod_725 <- mkDebugOperation(mod_725_inner, "mod_725");
    Operation_IFC mod_726_inner <- mkRepeatStatic(8);
    Operation_IFC mod_726 <- mkDebugOperation(mod_726_inner, "mod_726");
    Operation_IFC mod_727_inner <- mkFlatten(1);
    Operation_IFC mod_727 <- mkDebugOperation(mod_727_inner, "mod_727");
    Operation_IFC mod_728_inner <- mkFlatten(0);
    Operation_IFC mod_728 <- mkDebugOperation(mod_728_inner, "mod_728");
    PMU_IFC mod_729_bufferize <- mkPMU(1);
    Operation_IFC mod_729_inner = mod_729_bufferize.operation;
    Operation_IFC mod_729 <- mkDebugOperation(mod_729_inner, "mod_729");
    Operation_IFC mod_730_inner <- mkRepeatStatic(16);
    Operation_IFC mod_730 <- mkDebugOperation(mod_730_inner, "mod_730");
    PMU_IFC mod_731_bufferize <- mkPMU(2);
    Operation_IFC mod_731_inner = mod_731_bufferize.operation;
    Operation_IFC mod_731 <- mkDebugOperation(mod_731_inner, "mod_731");
    Operation_IFC mod_732_inner <- mkRepeatStatic(8);
    Operation_IFC mod_732 <- mkDebugOperation(mod_732_inner, "mod_732");
    Operation_IFC mod_733_inner <- mkFlatten(1);
    Operation_IFC mod_733 <- mkDebugOperation(mod_733_inner, "mod_733");
    Operation_IFC mod_734_inner <- mkFlatten(0);
    Operation_IFC mod_734 <- mkDebugOperation(mod_734_inner, "mod_734");
    Operation_IFC mod_735_inner <- mkRepeatStatic(16);
    Operation_IFC mod_735 <- mkDebugOperation(mod_735_inner, "mod_735");
    Operation_IFC mod_736_inner <- mkRepeatStatic(2);
    Operation_IFC mod_736 <- mkDebugOperation(mod_736_inner, "mod_736");
    PMU_IFC mod_737_bufferize <- mkPMU(2);
    Operation_IFC mod_737_inner = mod_737_bufferize.operation;
    Operation_IFC mod_737 <- mkDebugOperation(mod_737_inner, "mod_737");
    rule rule_902;
        ChannelMessage t;
        t <- mod_706.get(0);
        mod_707.put(0, t);
    endrule
    rule rule_903;
        ChannelMessage t;
        t <- mod_737.get(1);
        mod_701.put(1, t);
    endrule
    rule rule_904;
        ChannelMessage t;
        t <- mod_699.get(0);
        mod_700.put(0, t);
    endrule
    rule rule_905;
        ChannelMessage t;
        t <- mod_721.get(0);
        mod_709.put(1, t);
    endrule
    rule rule_906;
        ChannelMessage t;
        t <- mod_710.get(0);
        mod_711.put(0, t);
    endrule
    rule rule_907;
        ChannelMessage t;
        t <- mod_700.get(0);
        mod_701.put(0, t);
    endrule
    rule rule_908;
        ChannelMessage t;
        t <- mod_719.get(0);
        mod_717.put(0, t);
    endrule
    rule rule_909;
        ChannelMessage t;
        t <- mod_701.get(1);
        mod_702.put(0, t);
    endrule
    rule rule_910;
        ChannelMessage t;
        t <- mod_736.get(0);
        mod_703.put(1, t);
    endrule
    rule rule_911;
        ChannelMessage t;
        t <- mod_705.get(0);
        mod_735.put(0, t);
    endrule
    rule rule_912;
        ChannelMessage t;
        t <- mod_731.get(1);
        mod_706.put(1, t);
    endrule
    rule rule_913;
        ChannelMessage t;
        t <- mod_709.get(0);
        mod_721.put(0, t);
    endrule
    rule rule_914;
        ChannelMessage t;
        t <- mod_717.get(1);
        mod_710.put(1, t);
    endrule
    rule rule_915;
        ChannelMessage t;
        t <- mod_713.get(1);
        mod_714.put(1, t);
    endrule
    rule rule_916;
        ChannelMessage t;
        t <- mod_720.get(0);
        mod_719.put(0, t);
    endrule
    rule rule_917;
        ChannelMessage t;
        t <- mod_737.get(0);
        mod_737.put(1, t);
    endrule
    rule rule_918;
        ChannelMessage t;
        t <- mod_731.get(0);
        mod_732.put(0, t);
    endrule
    rule rule_919;
        ChannelMessage t;
        t <- mod_727.get(0);
        mod_725.put(0, t);
    endrule
    rule rule_920;
        ChannelMessage t;
        t <- mod_712.get(1);
        mod_713.put(0, t);
    endrule
    rule rule_921;
        ChannelMessage t;
        t <- mod_733.get(0);
        mod_731.put(0, t);
    endrule
    rule rule_922;
        ChannelMessage t;
        t <- mod_722.get(0);
        mod_708.put(1, t);
    endrule
    rule rule_923;
        ChannelMessage t;
        t <- mod_730.get(0);
        mod_729.put(1, t);
    endrule
    rule rule_924;
        ChannelMessage t;
        t <- mod_709.get(1);
        mod_710.put(0, t);
    endrule
    rule rule_925;
        ChannelMessage t;
        t <- mod_725.get(0);
        mod_726.put(0, t);
    endrule
    rule rule_926;
        ChannelMessage t;
        t <- mod_698.get(0);
        mod_699.put(0, t);
    endrule
    rule rule_927;
        ChannelMessage t;
        t <- mod_726.get(0);
        mod_725.put(1, t);
    endrule
    rule rule_928;
        ChannelMessage t;
        t <- mod_708.get(0);
        mod_709.put(0, t);
    endrule
    rule rule_929;
        ChannelMessage t;
        t <- mod_735.get(0);
        mod_705.put(1, t);
    endrule
    rule rule_930;
        ChannelMessage t;
        t <- mod_717.get(0);
        mod_718.put(0, t);
    endrule
    rule rule_931;
        ChannelMessage t;
        t <- mod_716.get(1);
        mod_712.put(1, t);
    endrule
    rule rule_932;
        ChannelMessage t;
        t <- mod_724.get(0);
        mod_723.put(0, t);
    endrule
    rule rule_933;
        ChannelMessage t;
        t <- mod_711.get(0);
        mod_712.put(0, t);
    endrule
    rule rule_934;
        ChannelMessage t;
        t <- mod_734.get(0);
        mod_733.put(0, t);
    endrule
    rule rule_935;
        ChannelMessage t;
        t <- mod_715.get(0);
        mod_715.put(1, t);
    endrule
    rule rule_936;
        ChannelMessage t;
        t <- mod_725.get(1);
        mod_724.put(1, t);
    endrule
    rule rule_937;
        ChannelMessage t;
        t <- mod_716.get(0);
        mod_716.put(1, t);
    endrule
    rule rule_938;
        ChannelMessage t;
        t <- mod_703.get(1);
        mod_704.put(0, t);
    endrule
    rule rule_939;
        ChannelMessage t;
        t <- mod_729.get(0);
        mod_730.put(0, t);
    endrule
    rule rule_940;
        ChannelMessage t;
        t <- mod_718.get(0);
        mod_717.put(1, t);
    endrule
    rule rule_941;
        ChannelMessage t;
        t <- mod_729.get(1);
        mod_724.put(0, t);
    endrule
    rule rule_942;
        ChannelMessage t;
        t <- mod_704.get(1);
        mod_705.put(0, t);
    endrule
    rule rule_943;
        ChannelMessage t;
        t <- mod_701.get(0);
        mod_737.put(0, t);
    endrule
    rule rule_944;
        ChannelMessage t;
        t <- mod_723.get(0);
        mod_722.put(0, t);
    endrule
    rule rule_945;
        ChannelMessage t;
        t <- mod_728.get(0);
        mod_727.put(0, t);
    endrule
    rule rule_946;
        ChannelMessage t;
        t <- mod_705.get(1);
        mod_706.put(0, t);
    endrule
    rule rule_947;
        ChannelMessage t;
        t <- mod_713.get(0);
        mod_715.put(0, t);
    endrule
    rule rule_948;
        ChannelMessage t;
        t <- mod_702.get(3);
        mod_703.put(0, t);
    endrule
    rule rule_949;
        ChannelMessage t;
        t <- mod_712.get(0);
        mod_716.put(0, t);
    endrule
    rule rule_950;
        ChannelMessage t;
        t <- mod_715.get(1);
        mod_713.put(1, t);
    endrule
    rule rule_951;
        ChannelMessage t;
        t <- mod_732.get(0);
        mod_731.put(1, t);
    endrule
    rule rule_952;
        ChannelMessage t;
        t <- mod_707.get(0);
        mod_708.put(0, t);
    endrule
    rule rule_953;
        ChannelMessage t;
        t <- mod_703.get(0);
        mod_736.put(0, t);
    endrule
    rule rule_954;
        ChannelMessage t;
        t <- mod_704.get(0);
        mod_729.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_698.put(0, t);
        end
        if (i == 1) begin
            mod_714.put(0, t);
        end
        if (i == 2) begin
            mod_720.put(0, t);
        end
        if (i == 3) begin
            mod_728.put(0, t);
        end
        if (i == 4) begin
            mod_734.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_702.get(0);
        end
        if (i == 2) begin
            t <- mod_702.get(1);
        end
        if (i == 0) begin
            t <- mod_702.get(2);
        end
        if (i == 1) begin
            t <- mod_714.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6052 (Operation_IFC);
    Operation_IFC mod_739_inner <- mkReshape(2, 64);
    Operation_IFC mod_739 <- mkDebugOperation(mod_739_inner, "mod_739");
    Operation_IFC mod_740_inner <- mkFlatten(1);
    Operation_IFC mod_740 <- mkDebugOperation(mod_740_inner, "mod_740");
    Operation_IFC mod_741_inner <- mkFlatten(2);
    Operation_IFC mod_741 <- mkDebugOperation(mod_741_inner, "mod_741");
    Operation_IFC mod_742_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_742 <- mkDebugOperation(mod_742_inner, "mod_742");
    Broadcast_IFC#(4) mod_743_inner <- mkBroadcast(4);
    Operation_IFC mod_743 <- mkDebugOperation(mod_743_inner.op, "mod_743");
    PMU_IFC mod_744_bufferize <- mkPMU(2);
    Operation_IFC mod_744_inner = mod_744_bufferize.operation;
    Operation_IFC mod_744 <- mkDebugOperation(mod_744_inner, "mod_744");
    Broadcast_IFC#(2) mod_745_inner <- mkBroadcast(2);
    Operation_IFC mod_745 <- mkDebugOperation(mod_745_inner.op, "mod_745");
    PMU_IFC mod_746_bufferize <- mkPMU(1);
    Operation_IFC mod_746_inner = mod_746_bufferize.operation;
    Operation_IFC mod_746 <- mkDebugOperation(mod_746_inner, "mod_746");
    Operation_IFC mod_747_inner <- mkBinaryMap(1138, matmul_t_tile);
    Operation_IFC mod_747 <- mkDebugOperation(mod_747_inner, "mod_747");
    Operation_IFC mod_748_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_748 <- mkDebugOperation(mod_748_inner, "mod_748");
    Operation_IFC mod_749_inner <- mkBinaryMap(1906, mul_tile);
    Operation_IFC mod_749 <- mkDebugOperation(mod_749_inner, "mod_749");
    PMU_IFC mod_750_bufferize <- mkPMU(1);
    Operation_IFC mod_750_inner = mod_750_bufferize.operation;
    Operation_IFC mod_750 <- mkDebugOperation(mod_750_inner, "mod_750");
    Operation_IFC mod_751_inner <- mkBinaryMap(2527, matmul_t_tile);
    Operation_IFC mod_751 <- mkDebugOperation(mod_751_inner, "mod_751");
    Operation_IFC mod_752_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_752 <- mkDebugOperation(mod_752_inner, "mod_752");
    Operation_IFC mod_753_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_753 <- mkDebugOperation(mod_753_inner, "mod_753");
    Operation_IFC mod_754_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_754 <- mkDebugOperation(mod_754_inner, "mod_754");
    Operation_IFC mod_755_inner <- mkBinaryMap(2805, mul_tile);
    Operation_IFC mod_755 <- mkDebugOperation(mod_755_inner, "mod_755");
    PMU_IFC mod_756_bufferize <- mkPMU(1);
    Operation_IFC mod_756_inner = mod_756_bufferize.operation;
    Operation_IFC mod_756 <- mkDebugOperation(mod_756_inner, "mod_756");
    PMU_IFC mod_757_bufferize <- mkPMU(2);
    Operation_IFC mod_757_inner = mod_757_bufferize.operation;
    Operation_IFC mod_757 <- mkDebugOperation(mod_757_inner, "mod_757");
    PMU_IFC mod_758_bufferize <- mkPMU(2);
    Operation_IFC mod_758_inner = mod_758_bufferize.operation;
    Operation_IFC mod_758 <- mkDebugOperation(mod_758_inner, "mod_758");
    Operation_IFC mod_759_inner <- mkRepeatStatic(8);
    Operation_IFC mod_759 <- mkDebugOperation(mod_759_inner, "mod_759");
    Operation_IFC mod_760_inner <- mkFlatten(1);
    Operation_IFC mod_760 <- mkDebugOperation(mod_760_inner, "mod_760");
    Operation_IFC mod_761_inner <- mkFlatten(0);
    Operation_IFC mod_761 <- mkDebugOperation(mod_761_inner, "mod_761");
    Operation_IFC mod_762_inner <- mkRepeatStatic(3);
    Operation_IFC mod_762 <- mkDebugOperation(mod_762_inner, "mod_762");
    Operation_IFC mod_763_inner <- mkUnaryMap(1778, silu_tile);
    Operation_IFC mod_763 <- mkDebugOperation(mod_763_inner, "mod_763");
    Operation_IFC mod_764_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_764 <- mkDebugOperation(mod_764_inner, "mod_764");
    Operation_IFC mod_765_inner <- mkBinaryMap(1650, matmul_t_tile);
    Operation_IFC mod_765 <- mkDebugOperation(mod_765_inner, "mod_765");
    PMU_IFC mod_766_bufferize <- mkPMU(2);
    Operation_IFC mod_766_inner = mod_766_bufferize.operation;
    Operation_IFC mod_766 <- mkDebugOperation(mod_766_inner, "mod_766");
    Operation_IFC mod_767_inner <- mkRepeatStatic(8);
    Operation_IFC mod_767 <- mkDebugOperation(mod_767_inner, "mod_767");
    Operation_IFC mod_768_inner <- mkFlatten(1);
    Operation_IFC mod_768 <- mkDebugOperation(mod_768_inner, "mod_768");
    Operation_IFC mod_769_inner <- mkFlatten(0);
    Operation_IFC mod_769 <- mkDebugOperation(mod_769_inner, "mod_769");
    PMU_IFC mod_770_bufferize <- mkPMU(1);
    Operation_IFC mod_770_inner = mod_770_bufferize.operation;
    Operation_IFC mod_770 <- mkDebugOperation(mod_770_inner, "mod_770");
    Operation_IFC mod_771_inner <- mkRepeatStatic(16);
    Operation_IFC mod_771 <- mkDebugOperation(mod_771_inner, "mod_771");
    PMU_IFC mod_772_bufferize <- mkPMU(2);
    Operation_IFC mod_772_inner = mod_772_bufferize.operation;
    Operation_IFC mod_772 <- mkDebugOperation(mod_772_inner, "mod_772");
    Operation_IFC mod_773_inner <- mkRepeatStatic(8);
    Operation_IFC mod_773 <- mkDebugOperation(mod_773_inner, "mod_773");
    Operation_IFC mod_774_inner <- mkFlatten(1);
    Operation_IFC mod_774 <- mkDebugOperation(mod_774_inner, "mod_774");
    Operation_IFC mod_775_inner <- mkFlatten(0);
    Operation_IFC mod_775 <- mkDebugOperation(mod_775_inner, "mod_775");
    Operation_IFC mod_776_inner <- mkRepeatStatic(16);
    Operation_IFC mod_776 <- mkDebugOperation(mod_776_inner, "mod_776");
    Operation_IFC mod_777_inner <- mkRepeatStatic(2);
    Operation_IFC mod_777 <- mkDebugOperation(mod_777_inner, "mod_777");
    PMU_IFC mod_778_bufferize <- mkPMU(2);
    Operation_IFC mod_778_inner = mod_778_bufferize.operation;
    Operation_IFC mod_778 <- mkDebugOperation(mod_778_inner, "mod_778");
    rule rule_955;
        ChannelMessage t;
        t <- mod_747.get(0);
        mod_748.put(0, t);
    endrule
    rule rule_956;
        ChannelMessage t;
        t <- mod_778.get(0);
        mod_778.put(1, t);
    endrule
    rule rule_957;
        ChannelMessage t;
        t <- mod_763.get(0);
        mod_749.put(1, t);
    endrule
    rule rule_958;
        ChannelMessage t;
        t <- mod_773.get(0);
        mod_772.put(1, t);
    endrule
    rule rule_959;
        ChannelMessage t;
        t <- mod_771.get(0);
        mod_770.put(1, t);
    endrule
    rule rule_960;
        ChannelMessage t;
        t <- mod_766.get(1);
        mod_765.put(1, t);
    endrule
    rule rule_961;
        ChannelMessage t;
        t <- mod_741.get(0);
        mod_742.put(0, t);
    endrule
    rule rule_962;
        ChannelMessage t;
        t <- mod_756.get(1);
        mod_754.put(1, t);
    endrule
    rule rule_963;
        ChannelMessage t;
        t <- mod_761.get(0);
        mod_760.put(0, t);
    endrule
    rule rule_964;
        ChannelMessage t;
        t <- mod_758.get(0);
        mod_759.put(0, t);
    endrule
    rule rule_965;
        ChannelMessage t;
        t <- mod_746.get(0);
        mod_776.put(0, t);
    endrule
    rule rule_966;
        ChannelMessage t;
        t <- mod_750.get(1);
        mod_751.put(0, t);
    endrule
    rule rule_967;
        ChannelMessage t;
        t <- mod_768.get(0);
        mod_766.put(0, t);
    endrule
    rule rule_968;
        ChannelMessage t;
        t <- mod_770.get(0);
        mod_771.put(0, t);
    endrule
    rule rule_969;
        ChannelMessage t;
        t <- mod_744.get(0);
        mod_777.put(0, t);
    endrule
    rule rule_970;
        ChannelMessage t;
        t <- mod_750.get(0);
        mod_762.put(0, t);
    endrule
    rule rule_971;
        ChannelMessage t;
        t <- mod_778.get(1);
        mod_742.put(1, t);
    endrule
    rule rule_972;
        ChannelMessage t;
        t <- mod_754.get(0);
        mod_756.put(0, t);
    endrule
    rule rule_973;
        ChannelMessage t;
        t <- mod_777.get(0);
        mod_744.put(1, t);
    endrule
    rule rule_974;
        ChannelMessage t;
        t <- mod_753.get(0);
        mod_757.put(0, t);
    endrule
    rule rule_975;
        ChannelMessage t;
        t <- mod_746.get(1);
        mod_747.put(0, t);
    endrule
    rule rule_976;
        ChannelMessage t;
        t <- mod_749.get(0);
        mod_750.put(0, t);
    endrule
    rule rule_977;
        ChannelMessage t;
        t <- mod_770.get(1);
        mod_765.put(0, t);
    endrule
    rule rule_978;
        ChannelMessage t;
        t <- mod_766.get(0);
        mod_767.put(0, t);
    endrule
    rule rule_979;
        ChannelMessage t;
        t <- mod_751.get(0);
        mod_752.put(0, t);
    endrule
    rule rule_980;
        ChannelMessage t;
        t <- mod_744.get(1);
        mod_745.put(0, t);
    endrule
    rule rule_981;
        ChannelMessage t;
        t <- mod_754.get(1);
        mod_755.put(1, t);
    endrule
    rule rule_982;
        ChannelMessage t;
        t <- mod_760.get(0);
        mod_758.put(0, t);
    endrule
    rule rule_983;
        ChannelMessage t;
        t <- mod_757.get(0);
        mod_757.put(1, t);
    endrule
    rule rule_984;
        ChannelMessage t;
        t <- mod_759.get(0);
        mod_758.put(1, t);
    endrule
    rule rule_985;
        ChannelMessage t;
        t <- mod_756.get(0);
        mod_756.put(1, t);
    endrule
    rule rule_986;
        ChannelMessage t;
        t <- mod_748.get(0);
        mod_749.put(0, t);
    endrule
    rule rule_987;
        ChannelMessage t;
        t <- mod_752.get(0);
        mod_753.put(0, t);
    endrule
    rule rule_988;
        ChannelMessage t;
        t <- mod_757.get(1);
        mod_753.put(1, t);
    endrule
    rule rule_989;
        ChannelMessage t;
        t <- mod_762.get(0);
        mod_750.put(1, t);
    endrule
    rule rule_990;
        ChannelMessage t;
        t <- mod_765.get(0);
        mod_764.put(0, t);
    endrule
    rule rule_991;
        ChannelMessage t;
        t <- mod_767.get(0);
        mod_766.put(1, t);
    endrule
    rule rule_992;
        ChannelMessage t;
        t <- mod_742.get(0);
        mod_778.put(0, t);
    endrule
    rule rule_993;
        ChannelMessage t;
        t <- mod_743.get(3);
        mod_744.put(0, t);
    endrule
    rule rule_994;
        ChannelMessage t;
        t <- mod_776.get(0);
        mod_746.put(1, t);
    endrule
    rule rule_995;
        ChannelMessage t;
        t <- mod_764.get(0);
        mod_763.put(0, t);
    endrule
    rule rule_996;
        ChannelMessage t;
        t <- mod_758.get(1);
        mod_751.put(1, t);
    endrule
    rule rule_997;
        ChannelMessage t;
        t <- mod_772.get(1);
        mod_747.put(1, t);
    endrule
    rule rule_998;
        ChannelMessage t;
        t <- mod_740.get(0);
        mod_741.put(0, t);
    endrule
    rule rule_999;
        ChannelMessage t;
        t <- mod_739.get(0);
        mod_740.put(0, t);
    endrule
    rule rule_1000;
        ChannelMessage t;
        t <- mod_742.get(1);
        mod_743.put(0, t);
    endrule
    rule rule_1001;
        ChannelMessage t;
        t <- mod_753.get(1);
        mod_754.put(0, t);
    endrule
    rule rule_1002;
        ChannelMessage t;
        t <- mod_769.get(0);
        mod_768.put(0, t);
    endrule
    rule rule_1003;
        ChannelMessage t;
        t <- mod_775.get(0);
        mod_774.put(0, t);
    endrule
    rule rule_1004;
        ChannelMessage t;
        t <- mod_745.get(0);
        mod_770.put(0, t);
    endrule
    rule rule_1005;
        ChannelMessage t;
        t <- mod_745.get(1);
        mod_746.put(0, t);
    endrule
    rule rule_1006;
        ChannelMessage t;
        t <- mod_774.get(0);
        mod_772.put(0, t);
    endrule
    rule rule_1007;
        ChannelMessage t;
        t <- mod_772.get(0);
        mod_773.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_739.put(0, t);
        end
        if (i == 1) begin
            mod_755.put(0, t);
        end
        if (i == 2) begin
            mod_761.put(0, t);
        end
        if (i == 3) begin
            mod_769.put(0, t);
        end
        if (i == 4) begin
            mod_775.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 2) begin
            t <- mod_743.get(0);
        end
        if (i == 1) begin
            t <- mod_743.get(1);
        end
        if (i == 0) begin
            t <- mod_743.get(2);
        end
        if (i == 3) begin
            t <- mod_755.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6053 (Operation_IFC);
    Operation_IFC mod_780_inner <- mkReshape(2, 64);
    Operation_IFC mod_780 <- mkDebugOperation(mod_780_inner, "mod_780");
    Operation_IFC mod_781_inner <- mkFlatten(1);
    Operation_IFC mod_781 <- mkDebugOperation(mod_781_inner, "mod_781");
    Operation_IFC mod_782_inner <- mkFlatten(2);
    Operation_IFC mod_782 <- mkDebugOperation(mod_782_inner, "mod_782");
    Operation_IFC mod_783_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_783 <- mkDebugOperation(mod_783_inner, "mod_783");
    Broadcast_IFC#(4) mod_784_inner <- mkBroadcast(4);
    Operation_IFC mod_784 <- mkDebugOperation(mod_784_inner.op, "mod_784");
    PMU_IFC mod_785_bufferize <- mkPMU(2);
    Operation_IFC mod_785_inner = mod_785_bufferize.operation;
    Operation_IFC mod_785 <- mkDebugOperation(mod_785_inner, "mod_785");
    Broadcast_IFC#(2) mod_786_inner <- mkBroadcast(2);
    Operation_IFC mod_786 <- mkDebugOperation(mod_786_inner.op, "mod_786");
    PMU_IFC mod_787_bufferize <- mkPMU(1);
    Operation_IFC mod_787_inner = mod_787_bufferize.operation;
    Operation_IFC mod_787 <- mkDebugOperation(mod_787_inner, "mod_787");
    Operation_IFC mod_788_inner <- mkBinaryMap(1137, matmul_t_tile);
    Operation_IFC mod_788 <- mkDebugOperation(mod_788_inner, "mod_788");
    Operation_IFC mod_789_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_789 <- mkDebugOperation(mod_789_inner, "mod_789");
    Operation_IFC mod_790_inner <- mkBinaryMap(1905, mul_tile);
    Operation_IFC mod_790 <- mkDebugOperation(mod_790_inner, "mod_790");
    PMU_IFC mod_791_bufferize <- mkPMU(1);
    Operation_IFC mod_791_inner = mod_791_bufferize.operation;
    Operation_IFC mod_791 <- mkDebugOperation(mod_791_inner, "mod_791");
    Operation_IFC mod_792_inner <- mkBinaryMap(2525, matmul_t_tile);
    Operation_IFC mod_792 <- mkDebugOperation(mod_792_inner, "mod_792");
    Operation_IFC mod_793_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_793 <- mkDebugOperation(mod_793_inner, "mod_793");
    Operation_IFC mod_794_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_794 <- mkDebugOperation(mod_794_inner, "mod_794");
    Operation_IFC mod_795_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_795 <- mkDebugOperation(mod_795_inner, "mod_795");
    Operation_IFC mod_796_inner <- mkBinaryMap(2804, mul_tile);
    Operation_IFC mod_796 <- mkDebugOperation(mod_796_inner, "mod_796");
    PMU_IFC mod_797_bufferize <- mkPMU(1);
    Operation_IFC mod_797_inner = mod_797_bufferize.operation;
    Operation_IFC mod_797 <- mkDebugOperation(mod_797_inner, "mod_797");
    PMU_IFC mod_798_bufferize <- mkPMU(2);
    Operation_IFC mod_798_inner = mod_798_bufferize.operation;
    Operation_IFC mod_798 <- mkDebugOperation(mod_798_inner, "mod_798");
    PMU_IFC mod_799_bufferize <- mkPMU(2);
    Operation_IFC mod_799_inner = mod_799_bufferize.operation;
    Operation_IFC mod_799 <- mkDebugOperation(mod_799_inner, "mod_799");
    Operation_IFC mod_800_inner <- mkRepeatStatic(8);
    Operation_IFC mod_800 <- mkDebugOperation(mod_800_inner, "mod_800");
    Operation_IFC mod_801_inner <- mkFlatten(1);
    Operation_IFC mod_801 <- mkDebugOperation(mod_801_inner, "mod_801");
    Operation_IFC mod_802_inner <- mkFlatten(0);
    Operation_IFC mod_802 <- mkDebugOperation(mod_802_inner, "mod_802");
    Operation_IFC mod_803_inner <- mkRepeatStatic(3);
    Operation_IFC mod_803 <- mkDebugOperation(mod_803_inner, "mod_803");
    Operation_IFC mod_804_inner <- mkUnaryMap(1777, silu_tile);
    Operation_IFC mod_804 <- mkDebugOperation(mod_804_inner, "mod_804");
    Operation_IFC mod_805_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_805 <- mkDebugOperation(mod_805_inner, "mod_805");
    Operation_IFC mod_806_inner <- mkBinaryMap(1649, matmul_t_tile);
    Operation_IFC mod_806 <- mkDebugOperation(mod_806_inner, "mod_806");
    PMU_IFC mod_807_bufferize <- mkPMU(2);
    Operation_IFC mod_807_inner = mod_807_bufferize.operation;
    Operation_IFC mod_807 <- mkDebugOperation(mod_807_inner, "mod_807");
    Operation_IFC mod_808_inner <- mkRepeatStatic(8);
    Operation_IFC mod_808 <- mkDebugOperation(mod_808_inner, "mod_808");
    Operation_IFC mod_809_inner <- mkFlatten(1);
    Operation_IFC mod_809 <- mkDebugOperation(mod_809_inner, "mod_809");
    Operation_IFC mod_810_inner <- mkFlatten(0);
    Operation_IFC mod_810 <- mkDebugOperation(mod_810_inner, "mod_810");
    PMU_IFC mod_811_bufferize <- mkPMU(1);
    Operation_IFC mod_811_inner = mod_811_bufferize.operation;
    Operation_IFC mod_811 <- mkDebugOperation(mod_811_inner, "mod_811");
    Operation_IFC mod_812_inner <- mkRepeatStatic(16);
    Operation_IFC mod_812 <- mkDebugOperation(mod_812_inner, "mod_812");
    PMU_IFC mod_813_bufferize <- mkPMU(2);
    Operation_IFC mod_813_inner = mod_813_bufferize.operation;
    Operation_IFC mod_813 <- mkDebugOperation(mod_813_inner, "mod_813");
    Operation_IFC mod_814_inner <- mkRepeatStatic(8);
    Operation_IFC mod_814 <- mkDebugOperation(mod_814_inner, "mod_814");
    Operation_IFC mod_815_inner <- mkFlatten(1);
    Operation_IFC mod_815 <- mkDebugOperation(mod_815_inner, "mod_815");
    Operation_IFC mod_816_inner <- mkFlatten(0);
    Operation_IFC mod_816 <- mkDebugOperation(mod_816_inner, "mod_816");
    Operation_IFC mod_817_inner <- mkRepeatStatic(16);
    Operation_IFC mod_817 <- mkDebugOperation(mod_817_inner, "mod_817");
    Operation_IFC mod_818_inner <- mkRepeatStatic(2);
    Operation_IFC mod_818 <- mkDebugOperation(mod_818_inner, "mod_818");
    PMU_IFC mod_819_bufferize <- mkPMU(2);
    Operation_IFC mod_819_inner = mod_819_bufferize.operation;
    Operation_IFC mod_819 <- mkDebugOperation(mod_819_inner, "mod_819");
    rule rule_1008;
        ChannelMessage t;
        t <- mod_791.get(0);
        mod_803.put(0, t);
    endrule
    rule rule_1009;
        ChannelMessage t;
        t <- mod_819.get(1);
        mod_783.put(1, t);
    endrule
    rule rule_1010;
        ChannelMessage t;
        t <- mod_806.get(0);
        mod_805.put(0, t);
    endrule
    rule rule_1011;
        ChannelMessage t;
        t <- mod_817.get(0);
        mod_787.put(1, t);
    endrule
    rule rule_1012;
        ChannelMessage t;
        t <- mod_800.get(0);
        mod_799.put(1, t);
    endrule
    rule rule_1013;
        ChannelMessage t;
        t <- mod_804.get(0);
        mod_790.put(1, t);
    endrule
    rule rule_1014;
        ChannelMessage t;
        t <- mod_783.get(1);
        mod_784.put(0, t);
    endrule
    rule rule_1015;
        ChannelMessage t;
        t <- mod_790.get(0);
        mod_791.put(0, t);
    endrule
    rule rule_1016;
        ChannelMessage t;
        t <- mod_810.get(0);
        mod_809.put(0, t);
    endrule
    rule rule_1017;
        ChannelMessage t;
        t <- mod_794.get(0);
        mod_798.put(0, t);
    endrule
    rule rule_1018;
        ChannelMessage t;
        t <- mod_797.get(0);
        mod_797.put(1, t);
    endrule
    rule rule_1019;
        ChannelMessage t;
        t <- mod_785.get(0);
        mod_818.put(0, t);
    endrule
    rule rule_1020;
        ChannelMessage t;
        t <- mod_812.get(0);
        mod_811.put(1, t);
    endrule
    rule rule_1021;
        ChannelMessage t;
        t <- mod_802.get(0);
        mod_801.put(0, t);
    endrule
    rule rule_1022;
        ChannelMessage t;
        t <- mod_786.get(1);
        mod_787.put(0, t);
    endrule
    rule rule_1023;
        ChannelMessage t;
        t <- mod_815.get(0);
        mod_813.put(0, t);
    endrule
    rule rule_1024;
        ChannelMessage t;
        t <- mod_795.get(0);
        mod_797.put(0, t);
    endrule
    rule rule_1025;
        ChannelMessage t;
        t <- mod_784.get(3);
        mod_785.put(0, t);
    endrule
    rule rule_1026;
        ChannelMessage t;
        t <- mod_808.get(0);
        mod_807.put(1, t);
    endrule
    rule rule_1027;
        ChannelMessage t;
        t <- mod_782.get(0);
        mod_783.put(0, t);
    endrule
    rule rule_1028;
        ChannelMessage t;
        t <- mod_795.get(1);
        mod_796.put(1, t);
    endrule
    rule rule_1029;
        ChannelMessage t;
        t <- mod_805.get(0);
        mod_804.put(0, t);
    endrule
    rule rule_1030;
        ChannelMessage t;
        t <- mod_811.get(0);
        mod_812.put(0, t);
    endrule
    rule rule_1031;
        ChannelMessage t;
        t <- mod_794.get(1);
        mod_795.put(0, t);
    endrule
    rule rule_1032;
        ChannelMessage t;
        t <- mod_785.get(1);
        mod_786.put(0, t);
    endrule
    rule rule_1033;
        ChannelMessage t;
        t <- mod_813.get(1);
        mod_788.put(1, t);
    endrule
    rule rule_1034;
        ChannelMessage t;
        t <- mod_801.get(0);
        mod_799.put(0, t);
    endrule
    rule rule_1035;
        ChannelMessage t;
        t <- mod_814.get(0);
        mod_813.put(1, t);
    endrule
    rule rule_1036;
        ChannelMessage t;
        t <- mod_807.get(0);
        mod_808.put(0, t);
    endrule
    rule rule_1037;
        ChannelMessage t;
        t <- mod_780.get(0);
        mod_781.put(0, t);
    endrule
    rule rule_1038;
        ChannelMessage t;
        t <- mod_793.get(0);
        mod_794.put(0, t);
    endrule
    rule rule_1039;
        ChannelMessage t;
        t <- mod_787.get(0);
        mod_817.put(0, t);
    endrule
    rule rule_1040;
        ChannelMessage t;
        t <- mod_788.get(0);
        mod_789.put(0, t);
    endrule
    rule rule_1041;
        ChannelMessage t;
        t <- mod_807.get(1);
        mod_806.put(1, t);
    endrule
    rule rule_1042;
        ChannelMessage t;
        t <- mod_786.get(0);
        mod_811.put(0, t);
    endrule
    rule rule_1043;
        ChannelMessage t;
        t <- mod_783.get(0);
        mod_819.put(0, t);
    endrule
    rule rule_1044;
        ChannelMessage t;
        t <- mod_798.get(1);
        mod_794.put(1, t);
    endrule
    rule rule_1045;
        ChannelMessage t;
        t <- mod_799.get(0);
        mod_800.put(0, t);
    endrule
    rule rule_1046;
        ChannelMessage t;
        t <- mod_813.get(0);
        mod_814.put(0, t);
    endrule
    rule rule_1047;
        ChannelMessage t;
        t <- mod_787.get(1);
        mod_788.put(0, t);
    endrule
    rule rule_1048;
        ChannelMessage t;
        t <- mod_798.get(0);
        mod_798.put(1, t);
    endrule
    rule rule_1049;
        ChannelMessage t;
        t <- mod_789.get(0);
        mod_790.put(0, t);
    endrule
    rule rule_1050;
        ChannelMessage t;
        t <- mod_797.get(1);
        mod_795.put(1, t);
    endrule
    rule rule_1051;
        ChannelMessage t;
        t <- mod_816.get(0);
        mod_815.put(0, t);
    endrule
    rule rule_1052;
        ChannelMessage t;
        t <- mod_809.get(0);
        mod_807.put(0, t);
    endrule
    rule rule_1053;
        ChannelMessage t;
        t <- mod_818.get(0);
        mod_785.put(1, t);
    endrule
    rule rule_1054;
        ChannelMessage t;
        t <- mod_781.get(0);
        mod_782.put(0, t);
    endrule
    rule rule_1055;
        ChannelMessage t;
        t <- mod_792.get(0);
        mod_793.put(0, t);
    endrule
    rule rule_1056;
        ChannelMessage t;
        t <- mod_803.get(0);
        mod_791.put(1, t);
    endrule
    rule rule_1057;
        ChannelMessage t;
        t <- mod_819.get(0);
        mod_819.put(1, t);
    endrule
    rule rule_1058;
        ChannelMessage t;
        t <- mod_791.get(1);
        mod_792.put(0, t);
    endrule
    rule rule_1059;
        ChannelMessage t;
        t <- mod_811.get(1);
        mod_806.put(0, t);
    endrule
    rule rule_1060;
        ChannelMessage t;
        t <- mod_799.get(1);
        mod_792.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_780.put(0, t);
        end
        if (i == 1) begin
            mod_796.put(0, t);
        end
        if (i == 2) begin
            mod_802.put(0, t);
        end
        if (i == 3) begin
            mod_810.put(0, t);
        end
        if (i == 4) begin
            mod_816.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_784.get(0);
        end
        if (i == 1) begin
            t <- mod_784.get(1);
        end
        if (i == 2) begin
            t <- mod_784.get(2);
        end
        if (i == 3) begin
            t <- mod_796.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6054 (Operation_IFC);
    Operation_IFC mod_821_inner <- mkReshape(2, 64);
    Operation_IFC mod_821 <- mkDebugOperation(mod_821_inner, "mod_821");
    Operation_IFC mod_822_inner <- mkFlatten(1);
    Operation_IFC mod_822 <- mkDebugOperation(mod_822_inner, "mod_822");
    Operation_IFC mod_823_inner <- mkFlatten(2);
    Operation_IFC mod_823 <- mkDebugOperation(mod_823_inner, "mod_823");
    Operation_IFC mod_824_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_824 <- mkDebugOperation(mod_824_inner, "mod_824");
    Broadcast_IFC#(4) mod_825_inner <- mkBroadcast(4);
    Operation_IFC mod_825 <- mkDebugOperation(mod_825_inner.op, "mod_825");
    PMU_IFC mod_826_bufferize <- mkPMU(2);
    Operation_IFC mod_826_inner = mod_826_bufferize.operation;
    Operation_IFC mod_826 <- mkDebugOperation(mod_826_inner, "mod_826");
    Broadcast_IFC#(2) mod_827_inner <- mkBroadcast(2);
    Operation_IFC mod_827 <- mkDebugOperation(mod_827_inner.op, "mod_827");
    PMU_IFC mod_828_bufferize <- mkPMU(1);
    Operation_IFC mod_828_inner = mod_828_bufferize.operation;
    Operation_IFC mod_828 <- mkDebugOperation(mod_828_inner, "mod_828");
    Operation_IFC mod_829_inner <- mkBinaryMap(1136, matmul_t_tile);
    Operation_IFC mod_829 <- mkDebugOperation(mod_829_inner, "mod_829");
    Operation_IFC mod_830_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_830 <- mkDebugOperation(mod_830_inner, "mod_830");
    Operation_IFC mod_831_inner <- mkBinaryMap(1904, mul_tile);
    Operation_IFC mod_831 <- mkDebugOperation(mod_831_inner, "mod_831");
    PMU_IFC mod_832_bufferize <- mkPMU(1);
    Operation_IFC mod_832_inner = mod_832_bufferize.operation;
    Operation_IFC mod_832 <- mkDebugOperation(mod_832_inner, "mod_832");
    Operation_IFC mod_833_inner <- mkBinaryMap(2523, matmul_t_tile);
    Operation_IFC mod_833 <- mkDebugOperation(mod_833_inner, "mod_833");
    Operation_IFC mod_834_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_834 <- mkDebugOperation(mod_834_inner, "mod_834");
    Operation_IFC mod_835_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_835 <- mkDebugOperation(mod_835_inner, "mod_835");
    Operation_IFC mod_836_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_836 <- mkDebugOperation(mod_836_inner, "mod_836");
    Operation_IFC mod_837_inner <- mkBinaryMap(2803, mul_tile);
    Operation_IFC mod_837 <- mkDebugOperation(mod_837_inner, "mod_837");
    PMU_IFC mod_838_bufferize <- mkPMU(1);
    Operation_IFC mod_838_inner = mod_838_bufferize.operation;
    Operation_IFC mod_838 <- mkDebugOperation(mod_838_inner, "mod_838");
    PMU_IFC mod_839_bufferize <- mkPMU(2);
    Operation_IFC mod_839_inner = mod_839_bufferize.operation;
    Operation_IFC mod_839 <- mkDebugOperation(mod_839_inner, "mod_839");
    PMU_IFC mod_840_bufferize <- mkPMU(2);
    Operation_IFC mod_840_inner = mod_840_bufferize.operation;
    Operation_IFC mod_840 <- mkDebugOperation(mod_840_inner, "mod_840");
    Operation_IFC mod_841_inner <- mkRepeatStatic(8);
    Operation_IFC mod_841 <- mkDebugOperation(mod_841_inner, "mod_841");
    Operation_IFC mod_842_inner <- mkFlatten(1);
    Operation_IFC mod_842 <- mkDebugOperation(mod_842_inner, "mod_842");
    Operation_IFC mod_843_inner <- mkFlatten(0);
    Operation_IFC mod_843 <- mkDebugOperation(mod_843_inner, "mod_843");
    Operation_IFC mod_844_inner <- mkRepeatStatic(3);
    Operation_IFC mod_844 <- mkDebugOperation(mod_844_inner, "mod_844");
    Operation_IFC mod_845_inner <- mkUnaryMap(1776, silu_tile);
    Operation_IFC mod_845 <- mkDebugOperation(mod_845_inner, "mod_845");
    Operation_IFC mod_846_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_846 <- mkDebugOperation(mod_846_inner, "mod_846");
    Operation_IFC mod_847_inner <- mkBinaryMap(1648, matmul_t_tile);
    Operation_IFC mod_847 <- mkDebugOperation(mod_847_inner, "mod_847");
    PMU_IFC mod_848_bufferize <- mkPMU(2);
    Operation_IFC mod_848_inner = mod_848_bufferize.operation;
    Operation_IFC mod_848 <- mkDebugOperation(mod_848_inner, "mod_848");
    Operation_IFC mod_849_inner <- mkRepeatStatic(8);
    Operation_IFC mod_849 <- mkDebugOperation(mod_849_inner, "mod_849");
    Operation_IFC mod_850_inner <- mkFlatten(1);
    Operation_IFC mod_850 <- mkDebugOperation(mod_850_inner, "mod_850");
    Operation_IFC mod_851_inner <- mkFlatten(0);
    Operation_IFC mod_851 <- mkDebugOperation(mod_851_inner, "mod_851");
    PMU_IFC mod_852_bufferize <- mkPMU(1);
    Operation_IFC mod_852_inner = mod_852_bufferize.operation;
    Operation_IFC mod_852 <- mkDebugOperation(mod_852_inner, "mod_852");
    Operation_IFC mod_853_inner <- mkRepeatStatic(16);
    Operation_IFC mod_853 <- mkDebugOperation(mod_853_inner, "mod_853");
    PMU_IFC mod_854_bufferize <- mkPMU(2);
    Operation_IFC mod_854_inner = mod_854_bufferize.operation;
    Operation_IFC mod_854 <- mkDebugOperation(mod_854_inner, "mod_854");
    Operation_IFC mod_855_inner <- mkRepeatStatic(8);
    Operation_IFC mod_855 <- mkDebugOperation(mod_855_inner, "mod_855");
    Operation_IFC mod_856_inner <- mkFlatten(1);
    Operation_IFC mod_856 <- mkDebugOperation(mod_856_inner, "mod_856");
    Operation_IFC mod_857_inner <- mkFlatten(0);
    Operation_IFC mod_857 <- mkDebugOperation(mod_857_inner, "mod_857");
    Operation_IFC mod_858_inner <- mkRepeatStatic(16);
    Operation_IFC mod_858 <- mkDebugOperation(mod_858_inner, "mod_858");
    Operation_IFC mod_859_inner <- mkRepeatStatic(2);
    Operation_IFC mod_859 <- mkDebugOperation(mod_859_inner, "mod_859");
    PMU_IFC mod_860_bufferize <- mkPMU(2);
    Operation_IFC mod_860_inner = mod_860_bufferize.operation;
    Operation_IFC mod_860 <- mkDebugOperation(mod_860_inner, "mod_860");
    rule rule_1061;
        ChannelMessage t;
        t <- mod_854.get(1);
        mod_829.put(1, t);
    endrule
    rule rule_1062;
        ChannelMessage t;
        t <- mod_859.get(0);
        mod_826.put(1, t);
    endrule
    rule rule_1063;
        ChannelMessage t;
        t <- mod_860.get(0);
        mod_860.put(1, t);
    endrule
    rule rule_1064;
        ChannelMessage t;
        t <- mod_840.get(0);
        mod_841.put(0, t);
    endrule
    rule rule_1065;
        ChannelMessage t;
        t <- mod_826.get(1);
        mod_827.put(0, t);
    endrule
    rule rule_1066;
        ChannelMessage t;
        t <- mod_827.get(1);
        mod_828.put(0, t);
    endrule
    rule rule_1067;
        ChannelMessage t;
        t <- mod_833.get(0);
        mod_834.put(0, t);
    endrule
    rule rule_1068;
        ChannelMessage t;
        t <- mod_851.get(0);
        mod_850.put(0, t);
    endrule
    rule rule_1069;
        ChannelMessage t;
        t <- mod_842.get(0);
        mod_840.put(0, t);
    endrule
    rule rule_1070;
        ChannelMessage t;
        t <- mod_845.get(0);
        mod_831.put(1, t);
    endrule
    rule rule_1071;
        ChannelMessage t;
        t <- mod_824.get(0);
        mod_860.put(0, t);
    endrule
    rule rule_1072;
        ChannelMessage t;
        t <- mod_834.get(0);
        mod_835.put(0, t);
    endrule
    rule rule_1073;
        ChannelMessage t;
        t <- mod_843.get(0);
        mod_842.put(0, t);
    endrule
    rule rule_1074;
        ChannelMessage t;
        t <- mod_847.get(0);
        mod_846.put(0, t);
    endrule
    rule rule_1075;
        ChannelMessage t;
        t <- mod_853.get(0);
        mod_852.put(1, t);
    endrule
    rule rule_1076;
        ChannelMessage t;
        t <- mod_832.get(1);
        mod_833.put(0, t);
    endrule
    rule rule_1077;
        ChannelMessage t;
        t <- mod_822.get(0);
        mod_823.put(0, t);
    endrule
    rule rule_1078;
        ChannelMessage t;
        t <- mod_838.get(1);
        mod_836.put(1, t);
    endrule
    rule rule_1079;
        ChannelMessage t;
        t <- mod_850.get(0);
        mod_848.put(0, t);
    endrule
    rule rule_1080;
        ChannelMessage t;
        t <- mod_827.get(0);
        mod_852.put(0, t);
    endrule
    rule rule_1081;
        ChannelMessage t;
        t <- mod_849.get(0);
        mod_848.put(1, t);
    endrule
    rule rule_1082;
        ChannelMessage t;
        t <- mod_841.get(0);
        mod_840.put(1, t);
    endrule
    rule rule_1083;
        ChannelMessage t;
        t <- mod_832.get(0);
        mod_844.put(0, t);
    endrule
    rule rule_1084;
        ChannelMessage t;
        t <- mod_823.get(0);
        mod_824.put(0, t);
    endrule
    rule rule_1085;
        ChannelMessage t;
        t <- mod_856.get(0);
        mod_854.put(0, t);
    endrule
    rule rule_1086;
        ChannelMessage t;
        t <- mod_836.get(1);
        mod_837.put(1, t);
    endrule
    rule rule_1087;
        ChannelMessage t;
        t <- mod_821.get(0);
        mod_822.put(0, t);
    endrule
    rule rule_1088;
        ChannelMessage t;
        t <- mod_840.get(1);
        mod_833.put(1, t);
    endrule
    rule rule_1089;
        ChannelMessage t;
        t <- mod_860.get(1);
        mod_824.put(1, t);
    endrule
    rule rule_1090;
        ChannelMessage t;
        t <- mod_839.get(1);
        mod_835.put(1, t);
    endrule
    rule rule_1091;
        ChannelMessage t;
        t <- mod_830.get(0);
        mod_831.put(0, t);
    endrule
    rule rule_1092;
        ChannelMessage t;
        t <- mod_828.get(1);
        mod_829.put(0, t);
    endrule
    rule rule_1093;
        ChannelMessage t;
        t <- mod_835.get(1);
        mod_836.put(0, t);
    endrule
    rule rule_1094;
        ChannelMessage t;
        t <- mod_854.get(0);
        mod_855.put(0, t);
    endrule
    rule rule_1095;
        ChannelMessage t;
        t <- mod_825.get(3);
        mod_826.put(0, t);
    endrule
    rule rule_1096;
        ChannelMessage t;
        t <- mod_852.get(0);
        mod_853.put(0, t);
    endrule
    rule rule_1097;
        ChannelMessage t;
        t <- mod_848.get(1);
        mod_847.put(1, t);
    endrule
    rule rule_1098;
        ChannelMessage t;
        t <- mod_855.get(0);
        mod_854.put(1, t);
    endrule
    rule rule_1099;
        ChannelMessage t;
        t <- mod_824.get(1);
        mod_825.put(0, t);
    endrule
    rule rule_1100;
        ChannelMessage t;
        t <- mod_829.get(0);
        mod_830.put(0, t);
    endrule
    rule rule_1101;
        ChannelMessage t;
        t <- mod_846.get(0);
        mod_845.put(0, t);
    endrule
    rule rule_1102;
        ChannelMessage t;
        t <- mod_848.get(0);
        mod_849.put(0, t);
    endrule
    rule rule_1103;
        ChannelMessage t;
        t <- mod_838.get(0);
        mod_838.put(1, t);
    endrule
    rule rule_1104;
        ChannelMessage t;
        t <- mod_836.get(0);
        mod_838.put(0, t);
    endrule
    rule rule_1105;
        ChannelMessage t;
        t <- mod_844.get(0);
        mod_832.put(1, t);
    endrule
    rule rule_1106;
        ChannelMessage t;
        t <- mod_831.get(0);
        mod_832.put(0, t);
    endrule
    rule rule_1107;
        ChannelMessage t;
        t <- mod_835.get(0);
        mod_839.put(0, t);
    endrule
    rule rule_1108;
        ChannelMessage t;
        t <- mod_839.get(0);
        mod_839.put(1, t);
    endrule
    rule rule_1109;
        ChannelMessage t;
        t <- mod_857.get(0);
        mod_856.put(0, t);
    endrule
    rule rule_1110;
        ChannelMessage t;
        t <- mod_858.get(0);
        mod_828.put(1, t);
    endrule
    rule rule_1111;
        ChannelMessage t;
        t <- mod_852.get(1);
        mod_847.put(0, t);
    endrule
    rule rule_1112;
        ChannelMessage t;
        t <- mod_828.get(0);
        mod_858.put(0, t);
    endrule
    rule rule_1113;
        ChannelMessage t;
        t <- mod_826.get(0);
        mod_859.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_821.put(0, t);
        end
        if (i == 1) begin
            mod_837.put(0, t);
        end
        if (i == 2) begin
            mod_843.put(0, t);
        end
        if (i == 3) begin
            mod_851.put(0, t);
        end
        if (i == 4) begin
            mod_857.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_825.get(0);
        end
        if (i == 1) begin
            t <- mod_825.get(1);
        end
        if (i == 3) begin
            t <- mod_825.get(2);
        end
        if (i == 2) begin
            t <- mod_837.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6055 (Operation_IFC);
    Operation_IFC mod_862_inner <- mkReshape(2, 64);
    Operation_IFC mod_862 <- mkDebugOperation(mod_862_inner, "mod_862");
    Operation_IFC mod_863_inner <- mkFlatten(1);
    Operation_IFC mod_863 <- mkDebugOperation(mod_863_inner, "mod_863");
    Operation_IFC mod_864_inner <- mkFlatten(2);
    Operation_IFC mod_864 <- mkDebugOperation(mod_864_inner, "mod_864");
    Operation_IFC mod_865_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_865 <- mkDebugOperation(mod_865_inner, "mod_865");
    Broadcast_IFC#(4) mod_866_inner <- mkBroadcast(4);
    Operation_IFC mod_866 <- mkDebugOperation(mod_866_inner.op, "mod_866");
    PMU_IFC mod_867_bufferize <- mkPMU(2);
    Operation_IFC mod_867_inner = mod_867_bufferize.operation;
    Operation_IFC mod_867 <- mkDebugOperation(mod_867_inner, "mod_867");
    Broadcast_IFC#(2) mod_868_inner <- mkBroadcast(2);
    Operation_IFC mod_868 <- mkDebugOperation(mod_868_inner.op, "mod_868");
    PMU_IFC mod_869_bufferize <- mkPMU(1);
    Operation_IFC mod_869_inner = mod_869_bufferize.operation;
    Operation_IFC mod_869 <- mkDebugOperation(mod_869_inner, "mod_869");
    Operation_IFC mod_870_inner <- mkBinaryMap(1135, matmul_t_tile);
    Operation_IFC mod_870 <- mkDebugOperation(mod_870_inner, "mod_870");
    Operation_IFC mod_871_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_871 <- mkDebugOperation(mod_871_inner, "mod_871");
    Operation_IFC mod_872_inner <- mkBinaryMap(1903, mul_tile);
    Operation_IFC mod_872 <- mkDebugOperation(mod_872_inner, "mod_872");
    PMU_IFC mod_873_bufferize <- mkPMU(1);
    Operation_IFC mod_873_inner = mod_873_bufferize.operation;
    Operation_IFC mod_873 <- mkDebugOperation(mod_873_inner, "mod_873");
    Operation_IFC mod_874_inner <- mkBinaryMap(2521, matmul_t_tile);
    Operation_IFC mod_874 <- mkDebugOperation(mod_874_inner, "mod_874");
    Operation_IFC mod_875_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_875 <- mkDebugOperation(mod_875_inner, "mod_875");
    Operation_IFC mod_876_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_876 <- mkDebugOperation(mod_876_inner, "mod_876");
    Operation_IFC mod_877_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_877 <- mkDebugOperation(mod_877_inner, "mod_877");
    Operation_IFC mod_878_inner <- mkBinaryMap(2802, mul_tile);
    Operation_IFC mod_878 <- mkDebugOperation(mod_878_inner, "mod_878");
    PMU_IFC mod_879_bufferize <- mkPMU(1);
    Operation_IFC mod_879_inner = mod_879_bufferize.operation;
    Operation_IFC mod_879 <- mkDebugOperation(mod_879_inner, "mod_879");
    PMU_IFC mod_880_bufferize <- mkPMU(2);
    Operation_IFC mod_880_inner = mod_880_bufferize.operation;
    Operation_IFC mod_880 <- mkDebugOperation(mod_880_inner, "mod_880");
    PMU_IFC mod_881_bufferize <- mkPMU(2);
    Operation_IFC mod_881_inner = mod_881_bufferize.operation;
    Operation_IFC mod_881 <- mkDebugOperation(mod_881_inner, "mod_881");
    Operation_IFC mod_882_inner <- mkRepeatStatic(8);
    Operation_IFC mod_882 <- mkDebugOperation(mod_882_inner, "mod_882");
    Operation_IFC mod_883_inner <- mkFlatten(1);
    Operation_IFC mod_883 <- mkDebugOperation(mod_883_inner, "mod_883");
    Operation_IFC mod_884_inner <- mkFlatten(0);
    Operation_IFC mod_884 <- mkDebugOperation(mod_884_inner, "mod_884");
    Operation_IFC mod_885_inner <- mkRepeatStatic(3);
    Operation_IFC mod_885 <- mkDebugOperation(mod_885_inner, "mod_885");
    Operation_IFC mod_886_inner <- mkUnaryMap(1775, silu_tile);
    Operation_IFC mod_886 <- mkDebugOperation(mod_886_inner, "mod_886");
    Operation_IFC mod_887_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_887 <- mkDebugOperation(mod_887_inner, "mod_887");
    Operation_IFC mod_888_inner <- mkBinaryMap(1647, matmul_t_tile);
    Operation_IFC mod_888 <- mkDebugOperation(mod_888_inner, "mod_888");
    PMU_IFC mod_889_bufferize <- mkPMU(2);
    Operation_IFC mod_889_inner = mod_889_bufferize.operation;
    Operation_IFC mod_889 <- mkDebugOperation(mod_889_inner, "mod_889");
    Operation_IFC mod_890_inner <- mkRepeatStatic(8);
    Operation_IFC mod_890 <- mkDebugOperation(mod_890_inner, "mod_890");
    Operation_IFC mod_891_inner <- mkFlatten(1);
    Operation_IFC mod_891 <- mkDebugOperation(mod_891_inner, "mod_891");
    Operation_IFC mod_892_inner <- mkFlatten(0);
    Operation_IFC mod_892 <- mkDebugOperation(mod_892_inner, "mod_892");
    PMU_IFC mod_893_bufferize <- mkPMU(1);
    Operation_IFC mod_893_inner = mod_893_bufferize.operation;
    Operation_IFC mod_893 <- mkDebugOperation(mod_893_inner, "mod_893");
    Operation_IFC mod_894_inner <- mkRepeatStatic(16);
    Operation_IFC mod_894 <- mkDebugOperation(mod_894_inner, "mod_894");
    PMU_IFC mod_895_bufferize <- mkPMU(2);
    Operation_IFC mod_895_inner = mod_895_bufferize.operation;
    Operation_IFC mod_895 <- mkDebugOperation(mod_895_inner, "mod_895");
    Operation_IFC mod_896_inner <- mkRepeatStatic(8);
    Operation_IFC mod_896 <- mkDebugOperation(mod_896_inner, "mod_896");
    Operation_IFC mod_897_inner <- mkFlatten(1);
    Operation_IFC mod_897 <- mkDebugOperation(mod_897_inner, "mod_897");
    Operation_IFC mod_898_inner <- mkFlatten(0);
    Operation_IFC mod_898 <- mkDebugOperation(mod_898_inner, "mod_898");
    Operation_IFC mod_899_inner <- mkRepeatStatic(16);
    Operation_IFC mod_899 <- mkDebugOperation(mod_899_inner, "mod_899");
    Operation_IFC mod_900_inner <- mkRepeatStatic(2);
    Operation_IFC mod_900 <- mkDebugOperation(mod_900_inner, "mod_900");
    PMU_IFC mod_901_bufferize <- mkPMU(2);
    Operation_IFC mod_901_inner = mod_901_bufferize.operation;
    Operation_IFC mod_901 <- mkDebugOperation(mod_901_inner, "mod_901");
    rule rule_1114;
        ChannelMessage t;
        t <- mod_868.get(0);
        mod_893.put(0, t);
    endrule
    rule rule_1115;
        ChannelMessage t;
        t <- mod_877.get(1);
        mod_878.put(1, t);
    endrule
    rule rule_1116;
        ChannelMessage t;
        t <- mod_889.get(1);
        mod_888.put(1, t);
    endrule
    rule rule_1117;
        ChannelMessage t;
        t <- mod_872.get(0);
        mod_873.put(0, t);
    endrule
    rule rule_1118;
        ChannelMessage t;
        t <- mod_871.get(0);
        mod_872.put(0, t);
    endrule
    rule rule_1119;
        ChannelMessage t;
        t <- mod_869.get(1);
        mod_870.put(0, t);
    endrule
    rule rule_1120;
        ChannelMessage t;
        t <- mod_882.get(0);
        mod_881.put(1, t);
    endrule
    rule rule_1121;
        ChannelMessage t;
        t <- mod_885.get(0);
        mod_873.put(1, t);
    endrule
    rule rule_1122;
        ChannelMessage t;
        t <- mod_890.get(0);
        mod_889.put(1, t);
    endrule
    rule rule_1123;
        ChannelMessage t;
        t <- mod_876.get(0);
        mod_880.put(0, t);
    endrule
    rule rule_1124;
        ChannelMessage t;
        t <- mod_862.get(0);
        mod_863.put(0, t);
    endrule
    rule rule_1125;
        ChannelMessage t;
        t <- mod_894.get(0);
        mod_893.put(1, t);
    endrule
    rule rule_1126;
        ChannelMessage t;
        t <- mod_887.get(0);
        mod_886.put(0, t);
    endrule
    rule rule_1127;
        ChannelMessage t;
        t <- mod_883.get(0);
        mod_881.put(0, t);
    endrule
    rule rule_1128;
        ChannelMessage t;
        t <- mod_873.get(1);
        mod_874.put(0, t);
    endrule
    rule rule_1129;
        ChannelMessage t;
        t <- mod_877.get(0);
        mod_879.put(0, t);
    endrule
    rule rule_1130;
        ChannelMessage t;
        t <- mod_864.get(0);
        mod_865.put(0, t);
    endrule
    rule rule_1131;
        ChannelMessage t;
        t <- mod_881.get(1);
        mod_874.put(1, t);
    endrule
    rule rule_1132;
        ChannelMessage t;
        t <- mod_895.get(1);
        mod_870.put(1, t);
    endrule
    rule rule_1133;
        ChannelMessage t;
        t <- mod_866.get(3);
        mod_867.put(0, t);
    endrule
    rule rule_1134;
        ChannelMessage t;
        t <- mod_889.get(0);
        mod_890.put(0, t);
    endrule
    rule rule_1135;
        ChannelMessage t;
        t <- mod_884.get(0);
        mod_883.put(0, t);
    endrule
    rule rule_1136;
        ChannelMessage t;
        t <- mod_865.get(1);
        mod_866.put(0, t);
    endrule
    rule rule_1137;
        ChannelMessage t;
        t <- mod_863.get(0);
        mod_864.put(0, t);
    endrule
    rule rule_1138;
        ChannelMessage t;
        t <- mod_870.get(0);
        mod_871.put(0, t);
    endrule
    rule rule_1139;
        ChannelMessage t;
        t <- mod_888.get(0);
        mod_887.put(0, t);
    endrule
    rule rule_1140;
        ChannelMessage t;
        t <- mod_891.get(0);
        mod_889.put(0, t);
    endrule
    rule rule_1141;
        ChannelMessage t;
        t <- mod_873.get(0);
        mod_885.put(0, t);
    endrule
    rule rule_1142;
        ChannelMessage t;
        t <- mod_900.get(0);
        mod_867.put(1, t);
    endrule
    rule rule_1143;
        ChannelMessage t;
        t <- mod_879.get(0);
        mod_879.put(1, t);
    endrule
    rule rule_1144;
        ChannelMessage t;
        t <- mod_867.get(1);
        mod_868.put(0, t);
    endrule
    rule rule_1145;
        ChannelMessage t;
        t <- mod_896.get(0);
        mod_895.put(1, t);
    endrule
    rule rule_1146;
        ChannelMessage t;
        t <- mod_869.get(0);
        mod_899.put(0, t);
    endrule
    rule rule_1147;
        ChannelMessage t;
        t <- mod_901.get(0);
        mod_901.put(1, t);
    endrule
    rule rule_1148;
        ChannelMessage t;
        t <- mod_867.get(0);
        mod_900.put(0, t);
    endrule
    rule rule_1149;
        ChannelMessage t;
        t <- mod_886.get(0);
        mod_872.put(1, t);
    endrule
    rule rule_1150;
        ChannelMessage t;
        t <- mod_897.get(0);
        mod_895.put(0, t);
    endrule
    rule rule_1151;
        ChannelMessage t;
        t <- mod_892.get(0);
        mod_891.put(0, t);
    endrule
    rule rule_1152;
        ChannelMessage t;
        t <- mod_865.get(0);
        mod_901.put(0, t);
    endrule
    rule rule_1153;
        ChannelMessage t;
        t <- mod_880.get(0);
        mod_880.put(1, t);
    endrule
    rule rule_1154;
        ChannelMessage t;
        t <- mod_880.get(1);
        mod_876.put(1, t);
    endrule
    rule rule_1155;
        ChannelMessage t;
        t <- mod_881.get(0);
        mod_882.put(0, t);
    endrule
    rule rule_1156;
        ChannelMessage t;
        t <- mod_895.get(0);
        mod_896.put(0, t);
    endrule
    rule rule_1157;
        ChannelMessage t;
        t <- mod_893.get(0);
        mod_894.put(0, t);
    endrule
    rule rule_1158;
        ChannelMessage t;
        t <- mod_874.get(0);
        mod_875.put(0, t);
    endrule
    rule rule_1159;
        ChannelMessage t;
        t <- mod_901.get(1);
        mod_865.put(1, t);
    endrule
    rule rule_1160;
        ChannelMessage t;
        t <- mod_876.get(1);
        mod_877.put(0, t);
    endrule
    rule rule_1161;
        ChannelMessage t;
        t <- mod_879.get(1);
        mod_877.put(1, t);
    endrule
    rule rule_1162;
        ChannelMessage t;
        t <- mod_899.get(0);
        mod_869.put(1, t);
    endrule
    rule rule_1163;
        ChannelMessage t;
        t <- mod_875.get(0);
        mod_876.put(0, t);
    endrule
    rule rule_1164;
        ChannelMessage t;
        t <- mod_898.get(0);
        mod_897.put(0, t);
    endrule
    rule rule_1165;
        ChannelMessage t;
        t <- mod_893.get(1);
        mod_888.put(0, t);
    endrule
    rule rule_1166;
        ChannelMessage t;
        t <- mod_868.get(1);
        mod_869.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_862.put(0, t);
        end
        if (i == 1) begin
            mod_878.put(0, t);
        end
        if (i == 2) begin
            mod_884.put(0, t);
        end
        if (i == 3) begin
            mod_892.put(0, t);
        end
        if (i == 4) begin
            mod_898.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_866.get(0);
        end
        if (i == 3) begin
            t <- mod_866.get(1);
        end
        if (i == 2) begin
            t <- mod_866.get(2);
        end
        if (i == 1) begin
            t <- mod_878.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6056 (Operation_IFC);
    Operation_IFC mod_903_inner <- mkReshape(2, 64);
    Operation_IFC mod_903 <- mkDebugOperation(mod_903_inner, "mod_903");
    Operation_IFC mod_904_inner <- mkFlatten(1);
    Operation_IFC mod_904 <- mkDebugOperation(mod_904_inner, "mod_904");
    Operation_IFC mod_905_inner <- mkFlatten(2);
    Operation_IFC mod_905 <- mkDebugOperation(mod_905_inner, "mod_905");
    Operation_IFC mod_906_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_906 <- mkDebugOperation(mod_906_inner, "mod_906");
    Broadcast_IFC#(4) mod_907_inner <- mkBroadcast(4);
    Operation_IFC mod_907 <- mkDebugOperation(mod_907_inner.op, "mod_907");
    PMU_IFC mod_908_bufferize <- mkPMU(2);
    Operation_IFC mod_908_inner = mod_908_bufferize.operation;
    Operation_IFC mod_908 <- mkDebugOperation(mod_908_inner, "mod_908");
    Broadcast_IFC#(2) mod_909_inner <- mkBroadcast(2);
    Operation_IFC mod_909 <- mkDebugOperation(mod_909_inner.op, "mod_909");
    PMU_IFC mod_910_bufferize <- mkPMU(1);
    Operation_IFC mod_910_inner = mod_910_bufferize.operation;
    Operation_IFC mod_910 <- mkDebugOperation(mod_910_inner, "mod_910");
    Operation_IFC mod_911_inner <- mkBinaryMap(1134, matmul_t_tile);
    Operation_IFC mod_911 <- mkDebugOperation(mod_911_inner, "mod_911");
    Operation_IFC mod_912_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_912 <- mkDebugOperation(mod_912_inner, "mod_912");
    Operation_IFC mod_913_inner <- mkBinaryMap(1902, mul_tile);
    Operation_IFC mod_913 <- mkDebugOperation(mod_913_inner, "mod_913");
    PMU_IFC mod_914_bufferize <- mkPMU(1);
    Operation_IFC mod_914_inner = mod_914_bufferize.operation;
    Operation_IFC mod_914 <- mkDebugOperation(mod_914_inner, "mod_914");
    Operation_IFC mod_915_inner <- mkBinaryMap(2519, matmul_t_tile);
    Operation_IFC mod_915 <- mkDebugOperation(mod_915_inner, "mod_915");
    Operation_IFC mod_916_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_916 <- mkDebugOperation(mod_916_inner, "mod_916");
    Operation_IFC mod_917_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_917 <- mkDebugOperation(mod_917_inner, "mod_917");
    Operation_IFC mod_918_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_918 <- mkDebugOperation(mod_918_inner, "mod_918");
    Operation_IFC mod_919_inner <- mkBinaryMap(2801, mul_tile);
    Operation_IFC mod_919 <- mkDebugOperation(mod_919_inner, "mod_919");
    PMU_IFC mod_920_bufferize <- mkPMU(1);
    Operation_IFC mod_920_inner = mod_920_bufferize.operation;
    Operation_IFC mod_920 <- mkDebugOperation(mod_920_inner, "mod_920");
    PMU_IFC mod_921_bufferize <- mkPMU(2);
    Operation_IFC mod_921_inner = mod_921_bufferize.operation;
    Operation_IFC mod_921 <- mkDebugOperation(mod_921_inner, "mod_921");
    PMU_IFC mod_922_bufferize <- mkPMU(2);
    Operation_IFC mod_922_inner = mod_922_bufferize.operation;
    Operation_IFC mod_922 <- mkDebugOperation(mod_922_inner, "mod_922");
    Operation_IFC mod_923_inner <- mkRepeatStatic(8);
    Operation_IFC mod_923 <- mkDebugOperation(mod_923_inner, "mod_923");
    Operation_IFC mod_924_inner <- mkFlatten(1);
    Operation_IFC mod_924 <- mkDebugOperation(mod_924_inner, "mod_924");
    Operation_IFC mod_925_inner <- mkFlatten(0);
    Operation_IFC mod_925 <- mkDebugOperation(mod_925_inner, "mod_925");
    Operation_IFC mod_926_inner <- mkRepeatStatic(3);
    Operation_IFC mod_926 <- mkDebugOperation(mod_926_inner, "mod_926");
    Operation_IFC mod_927_inner <- mkUnaryMap(1774, silu_tile);
    Operation_IFC mod_927 <- mkDebugOperation(mod_927_inner, "mod_927");
    Operation_IFC mod_928_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_928 <- mkDebugOperation(mod_928_inner, "mod_928");
    Operation_IFC mod_929_inner <- mkBinaryMap(1646, matmul_t_tile);
    Operation_IFC mod_929 <- mkDebugOperation(mod_929_inner, "mod_929");
    PMU_IFC mod_930_bufferize <- mkPMU(2);
    Operation_IFC mod_930_inner = mod_930_bufferize.operation;
    Operation_IFC mod_930 <- mkDebugOperation(mod_930_inner, "mod_930");
    Operation_IFC mod_931_inner <- mkRepeatStatic(8);
    Operation_IFC mod_931 <- mkDebugOperation(mod_931_inner, "mod_931");
    Operation_IFC mod_932_inner <- mkFlatten(1);
    Operation_IFC mod_932 <- mkDebugOperation(mod_932_inner, "mod_932");
    Operation_IFC mod_933_inner <- mkFlatten(0);
    Operation_IFC mod_933 <- mkDebugOperation(mod_933_inner, "mod_933");
    PMU_IFC mod_934_bufferize <- mkPMU(1);
    Operation_IFC mod_934_inner = mod_934_bufferize.operation;
    Operation_IFC mod_934 <- mkDebugOperation(mod_934_inner, "mod_934");
    Operation_IFC mod_935_inner <- mkRepeatStatic(16);
    Operation_IFC mod_935 <- mkDebugOperation(mod_935_inner, "mod_935");
    PMU_IFC mod_936_bufferize <- mkPMU(2);
    Operation_IFC mod_936_inner = mod_936_bufferize.operation;
    Operation_IFC mod_936 <- mkDebugOperation(mod_936_inner, "mod_936");
    Operation_IFC mod_937_inner <- mkRepeatStatic(8);
    Operation_IFC mod_937 <- mkDebugOperation(mod_937_inner, "mod_937");
    Operation_IFC mod_938_inner <- mkFlatten(1);
    Operation_IFC mod_938 <- mkDebugOperation(mod_938_inner, "mod_938");
    Operation_IFC mod_939_inner <- mkFlatten(0);
    Operation_IFC mod_939 <- mkDebugOperation(mod_939_inner, "mod_939");
    Operation_IFC mod_940_inner <- mkRepeatStatic(16);
    Operation_IFC mod_940 <- mkDebugOperation(mod_940_inner, "mod_940");
    Operation_IFC mod_941_inner <- mkRepeatStatic(2);
    Operation_IFC mod_941 <- mkDebugOperation(mod_941_inner, "mod_941");
    PMU_IFC mod_942_bufferize <- mkPMU(2);
    Operation_IFC mod_942_inner = mod_942_bufferize.operation;
    Operation_IFC mod_942 <- mkDebugOperation(mod_942_inner, "mod_942");
    rule rule_1167;
        ChannelMessage t;
        t <- mod_914.get(0);
        mod_926.put(0, t);
    endrule
    rule rule_1168;
        ChannelMessage t;
        t <- mod_909.get(0);
        mod_934.put(0, t);
    endrule
    rule rule_1169;
        ChannelMessage t;
        t <- mod_913.get(0);
        mod_914.put(0, t);
    endrule
    rule rule_1170;
        ChannelMessage t;
        t <- mod_918.get(1);
        mod_919.put(1, t);
    endrule
    rule rule_1171;
        ChannelMessage t;
        t <- mod_922.get(0);
        mod_923.put(0, t);
    endrule
    rule rule_1172;
        ChannelMessage t;
        t <- mod_930.get(0);
        mod_931.put(0, t);
    endrule
    rule rule_1173;
        ChannelMessage t;
        t <- mod_918.get(0);
        mod_920.put(0, t);
    endrule
    rule rule_1174;
        ChannelMessage t;
        t <- mod_936.get(1);
        mod_911.put(1, t);
    endrule
    rule rule_1175;
        ChannelMessage t;
        t <- mod_920.get(1);
        mod_918.put(1, t);
    endrule
    rule rule_1176;
        ChannelMessage t;
        t <- mod_921.get(1);
        mod_917.put(1, t);
    endrule
    rule rule_1177;
        ChannelMessage t;
        t <- mod_933.get(0);
        mod_932.put(0, t);
    endrule
    rule rule_1178;
        ChannelMessage t;
        t <- mod_907.get(3);
        mod_908.put(0, t);
    endrule
    rule rule_1179;
        ChannelMessage t;
        t <- mod_915.get(0);
        mod_916.put(0, t);
    endrule
    rule rule_1180;
        ChannelMessage t;
        t <- mod_923.get(0);
        mod_922.put(1, t);
    endrule
    rule rule_1181;
        ChannelMessage t;
        t <- mod_914.get(1);
        mod_915.put(0, t);
    endrule
    rule rule_1182;
        ChannelMessage t;
        t <- mod_937.get(0);
        mod_936.put(1, t);
    endrule
    rule rule_1183;
        ChannelMessage t;
        t <- mod_908.get(1);
        mod_909.put(0, t);
    endrule
    rule rule_1184;
        ChannelMessage t;
        t <- mod_931.get(0);
        mod_930.put(1, t);
    endrule
    rule rule_1185;
        ChannelMessage t;
        t <- mod_917.get(0);
        mod_921.put(0, t);
    endrule
    rule rule_1186;
        ChannelMessage t;
        t <- mod_921.get(0);
        mod_921.put(1, t);
    endrule
    rule rule_1187;
        ChannelMessage t;
        t <- mod_912.get(0);
        mod_913.put(0, t);
    endrule
    rule rule_1188;
        ChannelMessage t;
        t <- mod_909.get(1);
        mod_910.put(0, t);
    endrule
    rule rule_1189;
        ChannelMessage t;
        t <- mod_941.get(0);
        mod_908.put(1, t);
    endrule
    rule rule_1190;
        ChannelMessage t;
        t <- mod_911.get(0);
        mod_912.put(0, t);
    endrule
    rule rule_1191;
        ChannelMessage t;
        t <- mod_910.get(0);
        mod_940.put(0, t);
    endrule
    rule rule_1192;
        ChannelMessage t;
        t <- mod_934.get(1);
        mod_929.put(0, t);
    endrule
    rule rule_1193;
        ChannelMessage t;
        t <- mod_930.get(1);
        mod_929.put(1, t);
    endrule
    rule rule_1194;
        ChannelMessage t;
        t <- mod_922.get(1);
        mod_915.put(1, t);
    endrule
    rule rule_1195;
        ChannelMessage t;
        t <- mod_908.get(0);
        mod_941.put(0, t);
    endrule
    rule rule_1196;
        ChannelMessage t;
        t <- mod_932.get(0);
        mod_930.put(0, t);
    endrule
    rule rule_1197;
        ChannelMessage t;
        t <- mod_929.get(0);
        mod_928.put(0, t);
    endrule
    rule rule_1198;
        ChannelMessage t;
        t <- mod_942.get(0);
        mod_942.put(1, t);
    endrule
    rule rule_1199;
        ChannelMessage t;
        t <- mod_936.get(0);
        mod_937.put(0, t);
    endrule
    rule rule_1200;
        ChannelMessage t;
        t <- mod_938.get(0);
        mod_936.put(0, t);
    endrule
    rule rule_1201;
        ChannelMessage t;
        t <- mod_928.get(0);
        mod_927.put(0, t);
    endrule
    rule rule_1202;
        ChannelMessage t;
        t <- mod_924.get(0);
        mod_922.put(0, t);
    endrule
    rule rule_1203;
        ChannelMessage t;
        t <- mod_906.get(1);
        mod_907.put(0, t);
    endrule
    rule rule_1204;
        ChannelMessage t;
        t <- mod_925.get(0);
        mod_924.put(0, t);
    endrule
    rule rule_1205;
        ChannelMessage t;
        t <- mod_905.get(0);
        mod_906.put(0, t);
    endrule
    rule rule_1206;
        ChannelMessage t;
        t <- mod_942.get(1);
        mod_906.put(1, t);
    endrule
    rule rule_1207;
        ChannelMessage t;
        t <- mod_926.get(0);
        mod_914.put(1, t);
    endrule
    rule rule_1208;
        ChannelMessage t;
        t <- mod_910.get(1);
        mod_911.put(0, t);
    endrule
    rule rule_1209;
        ChannelMessage t;
        t <- mod_935.get(0);
        mod_934.put(1, t);
    endrule
    rule rule_1210;
        ChannelMessage t;
        t <- mod_903.get(0);
        mod_904.put(0, t);
    endrule
    rule rule_1211;
        ChannelMessage t;
        t <- mod_939.get(0);
        mod_938.put(0, t);
    endrule
    rule rule_1212;
        ChannelMessage t;
        t <- mod_927.get(0);
        mod_913.put(1, t);
    endrule
    rule rule_1213;
        ChannelMessage t;
        t <- mod_940.get(0);
        mod_910.put(1, t);
    endrule
    rule rule_1214;
        ChannelMessage t;
        t <- mod_934.get(0);
        mod_935.put(0, t);
    endrule
    rule rule_1215;
        ChannelMessage t;
        t <- mod_906.get(0);
        mod_942.put(0, t);
    endrule
    rule rule_1216;
        ChannelMessage t;
        t <- mod_917.get(1);
        mod_918.put(0, t);
    endrule
    rule rule_1217;
        ChannelMessage t;
        t <- mod_904.get(0);
        mod_905.put(0, t);
    endrule
    rule rule_1218;
        ChannelMessage t;
        t <- mod_916.get(0);
        mod_917.put(0, t);
    endrule
    rule rule_1219;
        ChannelMessage t;
        t <- mod_920.get(0);
        mod_920.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_903.put(0, t);
        end
        if (i == 1) begin
            mod_919.put(0, t);
        end
        if (i == 2) begin
            mod_925.put(0, t);
        end
        if (i == 3) begin
            mod_933.put(0, t);
        end
        if (i == 4) begin
            mod_939.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_907.get(0);
        end
        if (i == 2) begin
            t <- mod_907.get(1);
        end
        if (i == 3) begin
            t <- mod_907.get(2);
        end
        if (i == 1) begin
            t <- mod_919.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6057 (Operation_IFC);
    Operation_IFC mod_944_inner <- mkReshape(2, 64);
    Operation_IFC mod_944 <- mkDebugOperation(mod_944_inner, "mod_944");
    Operation_IFC mod_945_inner <- mkFlatten(1);
    Operation_IFC mod_945 <- mkDebugOperation(mod_945_inner, "mod_945");
    Operation_IFC mod_946_inner <- mkFlatten(2);
    Operation_IFC mod_946 <- mkDebugOperation(mod_946_inner, "mod_946");
    Operation_IFC mod_947_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_947 <- mkDebugOperation(mod_947_inner, "mod_947");
    Broadcast_IFC#(4) mod_948_inner <- mkBroadcast(4);
    Operation_IFC mod_948 <- mkDebugOperation(mod_948_inner.op, "mod_948");
    PMU_IFC mod_949_bufferize <- mkPMU(2);
    Operation_IFC mod_949_inner = mod_949_bufferize.operation;
    Operation_IFC mod_949 <- mkDebugOperation(mod_949_inner, "mod_949");
    Broadcast_IFC#(2) mod_950_inner <- mkBroadcast(2);
    Operation_IFC mod_950 <- mkDebugOperation(mod_950_inner.op, "mod_950");
    PMU_IFC mod_951_bufferize <- mkPMU(1);
    Operation_IFC mod_951_inner = mod_951_bufferize.operation;
    Operation_IFC mod_951 <- mkDebugOperation(mod_951_inner, "mod_951");
    Operation_IFC mod_952_inner <- mkBinaryMap(1133, matmul_t_tile);
    Operation_IFC mod_952 <- mkDebugOperation(mod_952_inner, "mod_952");
    Operation_IFC mod_953_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_953 <- mkDebugOperation(mod_953_inner, "mod_953");
    Operation_IFC mod_954_inner <- mkBinaryMap(1901, mul_tile);
    Operation_IFC mod_954 <- mkDebugOperation(mod_954_inner, "mod_954");
    PMU_IFC mod_955_bufferize <- mkPMU(1);
    Operation_IFC mod_955_inner = mod_955_bufferize.operation;
    Operation_IFC mod_955 <- mkDebugOperation(mod_955_inner, "mod_955");
    Operation_IFC mod_956_inner <- mkBinaryMap(2517, matmul_t_tile);
    Operation_IFC mod_956 <- mkDebugOperation(mod_956_inner, "mod_956");
    Operation_IFC mod_957_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_957 <- mkDebugOperation(mod_957_inner, "mod_957");
    Operation_IFC mod_958_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_958 <- mkDebugOperation(mod_958_inner, "mod_958");
    Operation_IFC mod_959_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_959 <- mkDebugOperation(mod_959_inner, "mod_959");
    Operation_IFC mod_960_inner <- mkBinaryMap(2800, mul_tile);
    Operation_IFC mod_960 <- mkDebugOperation(mod_960_inner, "mod_960");
    PMU_IFC mod_961_bufferize <- mkPMU(1);
    Operation_IFC mod_961_inner = mod_961_bufferize.operation;
    Operation_IFC mod_961 <- mkDebugOperation(mod_961_inner, "mod_961");
    PMU_IFC mod_962_bufferize <- mkPMU(2);
    Operation_IFC mod_962_inner = mod_962_bufferize.operation;
    Operation_IFC mod_962 <- mkDebugOperation(mod_962_inner, "mod_962");
    PMU_IFC mod_963_bufferize <- mkPMU(2);
    Operation_IFC mod_963_inner = mod_963_bufferize.operation;
    Operation_IFC mod_963 <- mkDebugOperation(mod_963_inner, "mod_963");
    Operation_IFC mod_964_inner <- mkRepeatStatic(8);
    Operation_IFC mod_964 <- mkDebugOperation(mod_964_inner, "mod_964");
    Operation_IFC mod_965_inner <- mkFlatten(1);
    Operation_IFC mod_965 <- mkDebugOperation(mod_965_inner, "mod_965");
    Operation_IFC mod_966_inner <- mkFlatten(0);
    Operation_IFC mod_966 <- mkDebugOperation(mod_966_inner, "mod_966");
    Operation_IFC mod_967_inner <- mkRepeatStatic(3);
    Operation_IFC mod_967 <- mkDebugOperation(mod_967_inner, "mod_967");
    Operation_IFC mod_968_inner <- mkUnaryMap(1773, silu_tile);
    Operation_IFC mod_968 <- mkDebugOperation(mod_968_inner, "mod_968");
    Operation_IFC mod_969_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_969 <- mkDebugOperation(mod_969_inner, "mod_969");
    Operation_IFC mod_970_inner <- mkBinaryMap(1645, matmul_t_tile);
    Operation_IFC mod_970 <- mkDebugOperation(mod_970_inner, "mod_970");
    PMU_IFC mod_971_bufferize <- mkPMU(2);
    Operation_IFC mod_971_inner = mod_971_bufferize.operation;
    Operation_IFC mod_971 <- mkDebugOperation(mod_971_inner, "mod_971");
    Operation_IFC mod_972_inner <- mkRepeatStatic(8);
    Operation_IFC mod_972 <- mkDebugOperation(mod_972_inner, "mod_972");
    Operation_IFC mod_973_inner <- mkFlatten(1);
    Operation_IFC mod_973 <- mkDebugOperation(mod_973_inner, "mod_973");
    Operation_IFC mod_974_inner <- mkFlatten(0);
    Operation_IFC mod_974 <- mkDebugOperation(mod_974_inner, "mod_974");
    PMU_IFC mod_975_bufferize <- mkPMU(1);
    Operation_IFC mod_975_inner = mod_975_bufferize.operation;
    Operation_IFC mod_975 <- mkDebugOperation(mod_975_inner, "mod_975");
    Operation_IFC mod_976_inner <- mkRepeatStatic(16);
    Operation_IFC mod_976 <- mkDebugOperation(mod_976_inner, "mod_976");
    PMU_IFC mod_977_bufferize <- mkPMU(2);
    Operation_IFC mod_977_inner = mod_977_bufferize.operation;
    Operation_IFC mod_977 <- mkDebugOperation(mod_977_inner, "mod_977");
    Operation_IFC mod_978_inner <- mkRepeatStatic(8);
    Operation_IFC mod_978 <- mkDebugOperation(mod_978_inner, "mod_978");
    Operation_IFC mod_979_inner <- mkFlatten(1);
    Operation_IFC mod_979 <- mkDebugOperation(mod_979_inner, "mod_979");
    Operation_IFC mod_980_inner <- mkFlatten(0);
    Operation_IFC mod_980 <- mkDebugOperation(mod_980_inner, "mod_980");
    Operation_IFC mod_981_inner <- mkRepeatStatic(16);
    Operation_IFC mod_981 <- mkDebugOperation(mod_981_inner, "mod_981");
    Operation_IFC mod_982_inner <- mkRepeatStatic(2);
    Operation_IFC mod_982 <- mkDebugOperation(mod_982_inner, "mod_982");
    PMU_IFC mod_983_bufferize <- mkPMU(2);
    Operation_IFC mod_983_inner = mod_983_bufferize.operation;
    Operation_IFC mod_983 <- mkDebugOperation(mod_983_inner, "mod_983");
    rule rule_1220;
        ChannelMessage t;
        t <- mod_975.get(0);
        mod_976.put(0, t);
    endrule
    rule rule_1221;
        ChannelMessage t;
        t <- mod_979.get(0);
        mod_977.put(0, t);
    endrule
    rule rule_1222;
        ChannelMessage t;
        t <- mod_980.get(0);
        mod_979.put(0, t);
    endrule
    rule rule_1223;
        ChannelMessage t;
        t <- mod_963.get(1);
        mod_956.put(1, t);
    endrule
    rule rule_1224;
        ChannelMessage t;
        t <- mod_961.get(0);
        mod_961.put(1, t);
    endrule
    rule rule_1225;
        ChannelMessage t;
        t <- mod_971.get(1);
        mod_970.put(1, t);
    endrule
    rule rule_1226;
        ChannelMessage t;
        t <- mod_961.get(1);
        mod_959.put(1, t);
    endrule
    rule rule_1227;
        ChannelMessage t;
        t <- mod_977.get(1);
        mod_952.put(1, t);
    endrule
    rule rule_1228;
        ChannelMessage t;
        t <- mod_945.get(0);
        mod_946.put(0, t);
    endrule
    rule rule_1229;
        ChannelMessage t;
        t <- mod_951.get(0);
        mod_981.put(0, t);
    endrule
    rule rule_1230;
        ChannelMessage t;
        t <- mod_944.get(0);
        mod_945.put(0, t);
    endrule
    rule rule_1231;
        ChannelMessage t;
        t <- mod_981.get(0);
        mod_951.put(1, t);
    endrule
    rule rule_1232;
        ChannelMessage t;
        t <- mod_951.get(1);
        mod_952.put(0, t);
    endrule
    rule rule_1233;
        ChannelMessage t;
        t <- mod_968.get(0);
        mod_954.put(1, t);
    endrule
    rule rule_1234;
        ChannelMessage t;
        t <- mod_974.get(0);
        mod_973.put(0, t);
    endrule
    rule rule_1235;
        ChannelMessage t;
        t <- mod_956.get(0);
        mod_957.put(0, t);
    endrule
    rule rule_1236;
        ChannelMessage t;
        t <- mod_978.get(0);
        mod_977.put(1, t);
    endrule
    rule rule_1237;
        ChannelMessage t;
        t <- mod_967.get(0);
        mod_955.put(1, t);
    endrule
    rule rule_1238;
        ChannelMessage t;
        t <- mod_947.get(1);
        mod_948.put(0, t);
    endrule
    rule rule_1239;
        ChannelMessage t;
        t <- mod_946.get(0);
        mod_947.put(0, t);
    endrule
    rule rule_1240;
        ChannelMessage t;
        t <- mod_962.get(0);
        mod_962.put(1, t);
    endrule
    rule rule_1241;
        ChannelMessage t;
        t <- mod_954.get(0);
        mod_955.put(0, t);
    endrule
    rule rule_1242;
        ChannelMessage t;
        t <- mod_948.get(3);
        mod_949.put(0, t);
    endrule
    rule rule_1243;
        ChannelMessage t;
        t <- mod_972.get(0);
        mod_971.put(1, t);
    endrule
    rule rule_1244;
        ChannelMessage t;
        t <- mod_958.get(0);
        mod_962.put(0, t);
    endrule
    rule rule_1245;
        ChannelMessage t;
        t <- mod_952.get(0);
        mod_953.put(0, t);
    endrule
    rule rule_1246;
        ChannelMessage t;
        t <- mod_949.get(0);
        mod_982.put(0, t);
    endrule
    rule rule_1247;
        ChannelMessage t;
        t <- mod_973.get(0);
        mod_971.put(0, t);
    endrule
    rule rule_1248;
        ChannelMessage t;
        t <- mod_950.get(1);
        mod_951.put(0, t);
    endrule
    rule rule_1249;
        ChannelMessage t;
        t <- mod_947.get(0);
        mod_983.put(0, t);
    endrule
    rule rule_1250;
        ChannelMessage t;
        t <- mod_958.get(1);
        mod_959.put(0, t);
    endrule
    rule rule_1251;
        ChannelMessage t;
        t <- mod_953.get(0);
        mod_954.put(0, t);
    endrule
    rule rule_1252;
        ChannelMessage t;
        t <- mod_955.get(1);
        mod_956.put(0, t);
    endrule
    rule rule_1253;
        ChannelMessage t;
        t <- mod_962.get(1);
        mod_958.put(1, t);
    endrule
    rule rule_1254;
        ChannelMessage t;
        t <- mod_966.get(0);
        mod_965.put(0, t);
    endrule
    rule rule_1255;
        ChannelMessage t;
        t <- mod_965.get(0);
        mod_963.put(0, t);
    endrule
    rule rule_1256;
        ChannelMessage t;
        t <- mod_971.get(0);
        mod_972.put(0, t);
    endrule
    rule rule_1257;
        ChannelMessage t;
        t <- mod_977.get(0);
        mod_978.put(0, t);
    endrule
    rule rule_1258;
        ChannelMessage t;
        t <- mod_983.get(1);
        mod_947.put(1, t);
    endrule
    rule rule_1259;
        ChannelMessage t;
        t <- mod_983.get(0);
        mod_983.put(1, t);
    endrule
    rule rule_1260;
        ChannelMessage t;
        t <- mod_982.get(0);
        mod_949.put(1, t);
    endrule
    rule rule_1261;
        ChannelMessage t;
        t <- mod_949.get(1);
        mod_950.put(0, t);
    endrule
    rule rule_1262;
        ChannelMessage t;
        t <- mod_959.get(1);
        mod_960.put(1, t);
    endrule
    rule rule_1263;
        ChannelMessage t;
        t <- mod_976.get(0);
        mod_975.put(1, t);
    endrule
    rule rule_1264;
        ChannelMessage t;
        t <- mod_950.get(0);
        mod_975.put(0, t);
    endrule
    rule rule_1265;
        ChannelMessage t;
        t <- mod_969.get(0);
        mod_968.put(0, t);
    endrule
    rule rule_1266;
        ChannelMessage t;
        t <- mod_975.get(1);
        mod_970.put(0, t);
    endrule
    rule rule_1267;
        ChannelMessage t;
        t <- mod_959.get(0);
        mod_961.put(0, t);
    endrule
    rule rule_1268;
        ChannelMessage t;
        t <- mod_964.get(0);
        mod_963.put(1, t);
    endrule
    rule rule_1269;
        ChannelMessage t;
        t <- mod_957.get(0);
        mod_958.put(0, t);
    endrule
    rule rule_1270;
        ChannelMessage t;
        t <- mod_955.get(0);
        mod_967.put(0, t);
    endrule
    rule rule_1271;
        ChannelMessage t;
        t <- mod_970.get(0);
        mod_969.put(0, t);
    endrule
    rule rule_1272;
        ChannelMessage t;
        t <- mod_963.get(0);
        mod_964.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_944.put(0, t);
        end
        if (i == 1) begin
            mod_960.put(0, t);
        end
        if (i == 2) begin
            mod_966.put(0, t);
        end
        if (i == 3) begin
            mod_974.put(0, t);
        end
        if (i == 4) begin
            mod_980.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_948.get(0);
        end
        if (i == 3) begin
            t <- mod_948.get(1);
        end
        if (i == 1) begin
            t <- mod_948.get(2);
        end
        if (i == 2) begin
            t <- mod_960.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6058 (Operation_IFC);
    Operation_IFC mod_985_inner <- mkReshape(2, 64);
    Operation_IFC mod_985 <- mkDebugOperation(mod_985_inner, "mod_985");
    Operation_IFC mod_986_inner <- mkFlatten(1);
    Operation_IFC mod_986 <- mkDebugOperation(mod_986_inner, "mod_986");
    Operation_IFC mod_987_inner <- mkFlatten(2);
    Operation_IFC mod_987 <- mkDebugOperation(mod_987_inner, "mod_987");
    Operation_IFC mod_988_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_988 <- mkDebugOperation(mod_988_inner, "mod_988");
    Broadcast_IFC#(4) mod_989_inner <- mkBroadcast(4);
    Operation_IFC mod_989 <- mkDebugOperation(mod_989_inner.op, "mod_989");
    PMU_IFC mod_990_bufferize <- mkPMU(2);
    Operation_IFC mod_990_inner = mod_990_bufferize.operation;
    Operation_IFC mod_990 <- mkDebugOperation(mod_990_inner, "mod_990");
    Broadcast_IFC#(2) mod_991_inner <- mkBroadcast(2);
    Operation_IFC mod_991 <- mkDebugOperation(mod_991_inner.op, "mod_991");
    PMU_IFC mod_992_bufferize <- mkPMU(1);
    Operation_IFC mod_992_inner = mod_992_bufferize.operation;
    Operation_IFC mod_992 <- mkDebugOperation(mod_992_inner, "mod_992");
    Operation_IFC mod_993_inner <- mkBinaryMap(1132, matmul_t_tile);
    Operation_IFC mod_993 <- mkDebugOperation(mod_993_inner, "mod_993");
    Operation_IFC mod_994_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_994 <- mkDebugOperation(mod_994_inner, "mod_994");
    Operation_IFC mod_995_inner <- mkBinaryMap(1900, mul_tile);
    Operation_IFC mod_995 <- mkDebugOperation(mod_995_inner, "mod_995");
    PMU_IFC mod_996_bufferize <- mkPMU(1);
    Operation_IFC mod_996_inner = mod_996_bufferize.operation;
    Operation_IFC mod_996 <- mkDebugOperation(mod_996_inner, "mod_996");
    Operation_IFC mod_997_inner <- mkBinaryMap(2515, matmul_t_tile);
    Operation_IFC mod_997 <- mkDebugOperation(mod_997_inner, "mod_997");
    Operation_IFC mod_998_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_998 <- mkDebugOperation(mod_998_inner, "mod_998");
    Operation_IFC mod_999_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_999 <- mkDebugOperation(mod_999_inner, "mod_999");
    Operation_IFC mod_1000_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1000 <- mkDebugOperation(mod_1000_inner, "mod_1000");
    Operation_IFC mod_1001_inner <- mkBinaryMap(2799, mul_tile);
    Operation_IFC mod_1001 <- mkDebugOperation(mod_1001_inner, "mod_1001");
    PMU_IFC mod_1002_bufferize <- mkPMU(1);
    Operation_IFC mod_1002_inner = mod_1002_bufferize.operation;
    Operation_IFC mod_1002 <- mkDebugOperation(mod_1002_inner, "mod_1002");
    PMU_IFC mod_1003_bufferize <- mkPMU(2);
    Operation_IFC mod_1003_inner = mod_1003_bufferize.operation;
    Operation_IFC mod_1003 <- mkDebugOperation(mod_1003_inner, "mod_1003");
    PMU_IFC mod_1004_bufferize <- mkPMU(2);
    Operation_IFC mod_1004_inner = mod_1004_bufferize.operation;
    Operation_IFC mod_1004 <- mkDebugOperation(mod_1004_inner, "mod_1004");
    Operation_IFC mod_1005_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1005 <- mkDebugOperation(mod_1005_inner, "mod_1005");
    Operation_IFC mod_1006_inner <- mkFlatten(1);
    Operation_IFC mod_1006 <- mkDebugOperation(mod_1006_inner, "mod_1006");
    Operation_IFC mod_1007_inner <- mkFlatten(0);
    Operation_IFC mod_1007 <- mkDebugOperation(mod_1007_inner, "mod_1007");
    Operation_IFC mod_1008_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1008 <- mkDebugOperation(mod_1008_inner, "mod_1008");
    Operation_IFC mod_1009_inner <- mkUnaryMap(1772, silu_tile);
    Operation_IFC mod_1009 <- mkDebugOperation(mod_1009_inner, "mod_1009");
    Operation_IFC mod_1010_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1010 <- mkDebugOperation(mod_1010_inner, "mod_1010");
    Operation_IFC mod_1011_inner <- mkBinaryMap(1644, matmul_t_tile);
    Operation_IFC mod_1011 <- mkDebugOperation(mod_1011_inner, "mod_1011");
    PMU_IFC mod_1012_bufferize <- mkPMU(2);
    Operation_IFC mod_1012_inner = mod_1012_bufferize.operation;
    Operation_IFC mod_1012 <- mkDebugOperation(mod_1012_inner, "mod_1012");
    Operation_IFC mod_1013_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1013 <- mkDebugOperation(mod_1013_inner, "mod_1013");
    Operation_IFC mod_1014_inner <- mkFlatten(1);
    Operation_IFC mod_1014 <- mkDebugOperation(mod_1014_inner, "mod_1014");
    Operation_IFC mod_1015_inner <- mkFlatten(0);
    Operation_IFC mod_1015 <- mkDebugOperation(mod_1015_inner, "mod_1015");
    PMU_IFC mod_1016_bufferize <- mkPMU(1);
    Operation_IFC mod_1016_inner = mod_1016_bufferize.operation;
    Operation_IFC mod_1016 <- mkDebugOperation(mod_1016_inner, "mod_1016");
    Operation_IFC mod_1017_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1017 <- mkDebugOperation(mod_1017_inner, "mod_1017");
    PMU_IFC mod_1018_bufferize <- mkPMU(2);
    Operation_IFC mod_1018_inner = mod_1018_bufferize.operation;
    Operation_IFC mod_1018 <- mkDebugOperation(mod_1018_inner, "mod_1018");
    Operation_IFC mod_1019_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1019 <- mkDebugOperation(mod_1019_inner, "mod_1019");
    Operation_IFC mod_1020_inner <- mkFlatten(1);
    Operation_IFC mod_1020 <- mkDebugOperation(mod_1020_inner, "mod_1020");
    Operation_IFC mod_1021_inner <- mkFlatten(0);
    Operation_IFC mod_1021 <- mkDebugOperation(mod_1021_inner, "mod_1021");
    Operation_IFC mod_1022_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1022 <- mkDebugOperation(mod_1022_inner, "mod_1022");
    Operation_IFC mod_1023_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1023 <- mkDebugOperation(mod_1023_inner, "mod_1023");
    PMU_IFC mod_1024_bufferize <- mkPMU(2);
    Operation_IFC mod_1024_inner = mod_1024_bufferize.operation;
    Operation_IFC mod_1024 <- mkDebugOperation(mod_1024_inner, "mod_1024");
    rule rule_1273;
        ChannelMessage t;
        t <- mod_1014.get(0);
        mod_1012.put(0, t);
    endrule
    rule rule_1274;
        ChannelMessage t;
        t <- mod_986.get(0);
        mod_987.put(0, t);
    endrule
    rule rule_1275;
        ChannelMessage t;
        t <- mod_1018.get(1);
        mod_993.put(1, t);
    endrule
    rule rule_1276;
        ChannelMessage t;
        t <- mod_989.get(3);
        mod_990.put(0, t);
    endrule
    rule rule_1277;
        ChannelMessage t;
        t <- mod_1012.get(1);
        mod_1011.put(1, t);
    endrule
    rule rule_1278;
        ChannelMessage t;
        t <- mod_1015.get(0);
        mod_1014.put(0, t);
    endrule
    rule rule_1279;
        ChannelMessage t;
        t <- mod_1004.get(0);
        mod_1005.put(0, t);
    endrule
    rule rule_1280;
        ChannelMessage t;
        t <- mod_996.get(0);
        mod_1008.put(0, t);
    endrule
    rule rule_1281;
        ChannelMessage t;
        t <- mod_1012.get(0);
        mod_1013.put(0, t);
    endrule
    rule rule_1282;
        ChannelMessage t;
        t <- mod_995.get(0);
        mod_996.put(0, t);
    endrule
    rule rule_1283;
        ChannelMessage t;
        t <- mod_1020.get(0);
        mod_1018.put(0, t);
    endrule
    rule rule_1284;
        ChannelMessage t;
        t <- mod_1000.get(0);
        mod_1002.put(0, t);
    endrule
    rule rule_1285;
        ChannelMessage t;
        t <- mod_1013.get(0);
        mod_1012.put(1, t);
    endrule
    rule rule_1286;
        ChannelMessage t;
        t <- mod_1005.get(0);
        mod_1004.put(1, t);
    endrule
    rule rule_1287;
        ChannelMessage t;
        t <- mod_1002.get(1);
        mod_1000.put(1, t);
    endrule
    rule rule_1288;
        ChannelMessage t;
        t <- mod_991.get(0);
        mod_1016.put(0, t);
    endrule
    rule rule_1289;
        ChannelMessage t;
        t <- mod_1019.get(0);
        mod_1018.put(1, t);
    endrule
    rule rule_1290;
        ChannelMessage t;
        t <- mod_1002.get(0);
        mod_1002.put(1, t);
    endrule
    rule rule_1291;
        ChannelMessage t;
        t <- mod_1004.get(1);
        mod_997.put(1, t);
    endrule
    rule rule_1292;
        ChannelMessage t;
        t <- mod_1017.get(0);
        mod_1016.put(1, t);
    endrule
    rule rule_1293;
        ChannelMessage t;
        t <- mod_1009.get(0);
        mod_995.put(1, t);
    endrule
    rule rule_1294;
        ChannelMessage t;
        t <- mod_1018.get(0);
        mod_1019.put(0, t);
    endrule
    rule rule_1295;
        ChannelMessage t;
        t <- mod_1008.get(0);
        mod_996.put(1, t);
    endrule
    rule rule_1296;
        ChannelMessage t;
        t <- mod_1003.get(0);
        mod_1003.put(1, t);
    endrule
    rule rule_1297;
        ChannelMessage t;
        t <- mod_988.get(0);
        mod_1024.put(0, t);
    endrule
    rule rule_1298;
        ChannelMessage t;
        t <- mod_987.get(0);
        mod_988.put(0, t);
    endrule
    rule rule_1299;
        ChannelMessage t;
        t <- mod_1000.get(1);
        mod_1001.put(1, t);
    endrule
    rule rule_1300;
        ChannelMessage t;
        t <- mod_1006.get(0);
        mod_1004.put(0, t);
    endrule
    rule rule_1301;
        ChannelMessage t;
        t <- mod_994.get(0);
        mod_995.put(0, t);
    endrule
    rule rule_1302;
        ChannelMessage t;
        t <- mod_999.get(0);
        mod_1003.put(0, t);
    endrule
    rule rule_1303;
        ChannelMessage t;
        t <- mod_998.get(0);
        mod_999.put(0, t);
    endrule
    rule rule_1304;
        ChannelMessage t;
        t <- mod_1024.get(1);
        mod_988.put(1, t);
    endrule
    rule rule_1305;
        ChannelMessage t;
        t <- mod_985.get(0);
        mod_986.put(0, t);
    endrule
    rule rule_1306;
        ChannelMessage t;
        t <- mod_996.get(1);
        mod_997.put(0, t);
    endrule
    rule rule_1307;
        ChannelMessage t;
        t <- mod_1011.get(0);
        mod_1010.put(0, t);
    endrule
    rule rule_1308;
        ChannelMessage t;
        t <- mod_1022.get(0);
        mod_992.put(1, t);
    endrule
    rule rule_1309;
        ChannelMessage t;
        t <- mod_992.get(0);
        mod_1022.put(0, t);
    endrule
    rule rule_1310;
        ChannelMessage t;
        t <- mod_993.get(0);
        mod_994.put(0, t);
    endrule
    rule rule_1311;
        ChannelMessage t;
        t <- mod_1003.get(1);
        mod_999.put(1, t);
    endrule
    rule rule_1312;
        ChannelMessage t;
        t <- mod_988.get(1);
        mod_989.put(0, t);
    endrule
    rule rule_1313;
        ChannelMessage t;
        t <- mod_997.get(0);
        mod_998.put(0, t);
    endrule
    rule rule_1314;
        ChannelMessage t;
        t <- mod_992.get(1);
        mod_993.put(0, t);
    endrule
    rule rule_1315;
        ChannelMessage t;
        t <- mod_1016.get(0);
        mod_1017.put(0, t);
    endrule
    rule rule_1316;
        ChannelMessage t;
        t <- mod_1016.get(1);
        mod_1011.put(0, t);
    endrule
    rule rule_1317;
        ChannelMessage t;
        t <- mod_999.get(1);
        mod_1000.put(0, t);
    endrule
    rule rule_1318;
        ChannelMessage t;
        t <- mod_1023.get(0);
        mod_990.put(1, t);
    endrule
    rule rule_1319;
        ChannelMessage t;
        t <- mod_991.get(1);
        mod_992.put(0, t);
    endrule
    rule rule_1320;
        ChannelMessage t;
        t <- mod_1007.get(0);
        mod_1006.put(0, t);
    endrule
    rule rule_1321;
        ChannelMessage t;
        t <- mod_990.get(1);
        mod_991.put(0, t);
    endrule
    rule rule_1322;
        ChannelMessage t;
        t <- mod_1021.get(0);
        mod_1020.put(0, t);
    endrule
    rule rule_1323;
        ChannelMessage t;
        t <- mod_1024.get(0);
        mod_1024.put(1, t);
    endrule
    rule rule_1324;
        ChannelMessage t;
        t <- mod_990.get(0);
        mod_1023.put(0, t);
    endrule
    rule rule_1325;
        ChannelMessage t;
        t <- mod_1010.get(0);
        mod_1009.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_985.put(0, t);
        end
        if (i == 1) begin
            mod_1001.put(0, t);
        end
        if (i == 2) begin
            mod_1007.put(0, t);
        end
        if (i == 3) begin
            mod_1015.put(0, t);
        end
        if (i == 4) begin
            mod_1021.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_989.get(0);
        end
        if (i == 2) begin
            t <- mod_989.get(1);
        end
        if (i == 0) begin
            t <- mod_989.get(2);
        end
        if (i == 3) begin
            t <- mod_1001.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6059 (Operation_IFC);
    Operation_IFC mod_1026_inner <- mkReshape(2, 64);
    Operation_IFC mod_1026 <- mkDebugOperation(mod_1026_inner, "mod_1026");
    Operation_IFC mod_1027_inner <- mkFlatten(1);
    Operation_IFC mod_1027 <- mkDebugOperation(mod_1027_inner, "mod_1027");
    Operation_IFC mod_1028_inner <- mkFlatten(2);
    Operation_IFC mod_1028 <- mkDebugOperation(mod_1028_inner, "mod_1028");
    Operation_IFC mod_1029_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1029 <- mkDebugOperation(mod_1029_inner, "mod_1029");
    Broadcast_IFC#(4) mod_1030_inner <- mkBroadcast(4);
    Operation_IFC mod_1030 <- mkDebugOperation(mod_1030_inner.op, "mod_1030");
    PMU_IFC mod_1031_bufferize <- mkPMU(2);
    Operation_IFC mod_1031_inner = mod_1031_bufferize.operation;
    Operation_IFC mod_1031 <- mkDebugOperation(mod_1031_inner, "mod_1031");
    Broadcast_IFC#(2) mod_1032_inner <- mkBroadcast(2);
    Operation_IFC mod_1032 <- mkDebugOperation(mod_1032_inner.op, "mod_1032");
    PMU_IFC mod_1033_bufferize <- mkPMU(1);
    Operation_IFC mod_1033_inner = mod_1033_bufferize.operation;
    Operation_IFC mod_1033 <- mkDebugOperation(mod_1033_inner, "mod_1033");
    Operation_IFC mod_1034_inner <- mkBinaryMap(1131, matmul_t_tile);
    Operation_IFC mod_1034 <- mkDebugOperation(mod_1034_inner, "mod_1034");
    Operation_IFC mod_1035_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1035 <- mkDebugOperation(mod_1035_inner, "mod_1035");
    Operation_IFC mod_1036_inner <- mkBinaryMap(1899, mul_tile);
    Operation_IFC mod_1036 <- mkDebugOperation(mod_1036_inner, "mod_1036");
    PMU_IFC mod_1037_bufferize <- mkPMU(1);
    Operation_IFC mod_1037_inner = mod_1037_bufferize.operation;
    Operation_IFC mod_1037 <- mkDebugOperation(mod_1037_inner, "mod_1037");
    Operation_IFC mod_1038_inner <- mkBinaryMap(2513, matmul_t_tile);
    Operation_IFC mod_1038 <- mkDebugOperation(mod_1038_inner, "mod_1038");
    Operation_IFC mod_1039_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1039 <- mkDebugOperation(mod_1039_inner, "mod_1039");
    Operation_IFC mod_1040_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1040 <- mkDebugOperation(mod_1040_inner, "mod_1040");
    Operation_IFC mod_1041_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1041 <- mkDebugOperation(mod_1041_inner, "mod_1041");
    Operation_IFC mod_1042_inner <- mkBinaryMap(2798, mul_tile);
    Operation_IFC mod_1042 <- mkDebugOperation(mod_1042_inner, "mod_1042");
    PMU_IFC mod_1043_bufferize <- mkPMU(1);
    Operation_IFC mod_1043_inner = mod_1043_bufferize.operation;
    Operation_IFC mod_1043 <- mkDebugOperation(mod_1043_inner, "mod_1043");
    PMU_IFC mod_1044_bufferize <- mkPMU(2);
    Operation_IFC mod_1044_inner = mod_1044_bufferize.operation;
    Operation_IFC mod_1044 <- mkDebugOperation(mod_1044_inner, "mod_1044");
    PMU_IFC mod_1045_bufferize <- mkPMU(2);
    Operation_IFC mod_1045_inner = mod_1045_bufferize.operation;
    Operation_IFC mod_1045 <- mkDebugOperation(mod_1045_inner, "mod_1045");
    Operation_IFC mod_1046_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1046 <- mkDebugOperation(mod_1046_inner, "mod_1046");
    Operation_IFC mod_1047_inner <- mkFlatten(1);
    Operation_IFC mod_1047 <- mkDebugOperation(mod_1047_inner, "mod_1047");
    Operation_IFC mod_1048_inner <- mkFlatten(0);
    Operation_IFC mod_1048 <- mkDebugOperation(mod_1048_inner, "mod_1048");
    Operation_IFC mod_1049_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1049 <- mkDebugOperation(mod_1049_inner, "mod_1049");
    Operation_IFC mod_1050_inner <- mkUnaryMap(1771, silu_tile);
    Operation_IFC mod_1050 <- mkDebugOperation(mod_1050_inner, "mod_1050");
    Operation_IFC mod_1051_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1051 <- mkDebugOperation(mod_1051_inner, "mod_1051");
    Operation_IFC mod_1052_inner <- mkBinaryMap(1643, matmul_t_tile);
    Operation_IFC mod_1052 <- mkDebugOperation(mod_1052_inner, "mod_1052");
    PMU_IFC mod_1053_bufferize <- mkPMU(2);
    Operation_IFC mod_1053_inner = mod_1053_bufferize.operation;
    Operation_IFC mod_1053 <- mkDebugOperation(mod_1053_inner, "mod_1053");
    Operation_IFC mod_1054_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1054 <- mkDebugOperation(mod_1054_inner, "mod_1054");
    Operation_IFC mod_1055_inner <- mkFlatten(1);
    Operation_IFC mod_1055 <- mkDebugOperation(mod_1055_inner, "mod_1055");
    Operation_IFC mod_1056_inner <- mkFlatten(0);
    Operation_IFC mod_1056 <- mkDebugOperation(mod_1056_inner, "mod_1056");
    PMU_IFC mod_1057_bufferize <- mkPMU(1);
    Operation_IFC mod_1057_inner = mod_1057_bufferize.operation;
    Operation_IFC mod_1057 <- mkDebugOperation(mod_1057_inner, "mod_1057");
    Operation_IFC mod_1058_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1058 <- mkDebugOperation(mod_1058_inner, "mod_1058");
    PMU_IFC mod_1059_bufferize <- mkPMU(2);
    Operation_IFC mod_1059_inner = mod_1059_bufferize.operation;
    Operation_IFC mod_1059 <- mkDebugOperation(mod_1059_inner, "mod_1059");
    Operation_IFC mod_1060_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1060 <- mkDebugOperation(mod_1060_inner, "mod_1060");
    Operation_IFC mod_1061_inner <- mkFlatten(1);
    Operation_IFC mod_1061 <- mkDebugOperation(mod_1061_inner, "mod_1061");
    Operation_IFC mod_1062_inner <- mkFlatten(0);
    Operation_IFC mod_1062 <- mkDebugOperation(mod_1062_inner, "mod_1062");
    Operation_IFC mod_1063_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1063 <- mkDebugOperation(mod_1063_inner, "mod_1063");
    Operation_IFC mod_1064_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1064 <- mkDebugOperation(mod_1064_inner, "mod_1064");
    PMU_IFC mod_1065_bufferize <- mkPMU(2);
    Operation_IFC mod_1065_inner = mod_1065_bufferize.operation;
    Operation_IFC mod_1065 <- mkDebugOperation(mod_1065_inner, "mod_1065");
    rule rule_1326;
        ChannelMessage t;
        t <- mod_1037.get(0);
        mod_1049.put(0, t);
    endrule
    rule rule_1327;
        ChannelMessage t;
        t <- mod_1062.get(0);
        mod_1061.put(0, t);
    endrule
    rule rule_1328;
        ChannelMessage t;
        t <- mod_1039.get(0);
        mod_1040.put(0, t);
    endrule
    rule rule_1329;
        ChannelMessage t;
        t <- mod_1032.get(0);
        mod_1057.put(0, t);
    endrule
    rule rule_1330;
        ChannelMessage t;
        t <- mod_1059.get(0);
        mod_1060.put(0, t);
    endrule
    rule rule_1331;
        ChannelMessage t;
        t <- mod_1064.get(0);
        mod_1031.put(1, t);
    endrule
    rule rule_1332;
        ChannelMessage t;
        t <- mod_1056.get(0);
        mod_1055.put(0, t);
    endrule
    rule rule_1333;
        ChannelMessage t;
        t <- mod_1065.get(0);
        mod_1065.put(1, t);
    endrule
    rule rule_1334;
        ChannelMessage t;
        t <- mod_1044.get(1);
        mod_1040.put(1, t);
    endrule
    rule rule_1335;
        ChannelMessage t;
        t <- mod_1038.get(0);
        mod_1039.put(0, t);
    endrule
    rule rule_1336;
        ChannelMessage t;
        t <- mod_1037.get(1);
        mod_1038.put(0, t);
    endrule
    rule rule_1337;
        ChannelMessage t;
        t <- mod_1050.get(0);
        mod_1036.put(1, t);
    endrule
    rule rule_1338;
        ChannelMessage t;
        t <- mod_1054.get(0);
        mod_1053.put(1, t);
    endrule
    rule rule_1339;
        ChannelMessage t;
        t <- mod_1030.get(3);
        mod_1031.put(0, t);
    endrule
    rule rule_1340;
        ChannelMessage t;
        t <- mod_1059.get(1);
        mod_1034.put(1, t);
    endrule
    rule rule_1341;
        ChannelMessage t;
        t <- mod_1052.get(0);
        mod_1051.put(0, t);
    endrule
    rule rule_1342;
        ChannelMessage t;
        t <- mod_1040.get(0);
        mod_1044.put(0, t);
    endrule
    rule rule_1343;
        ChannelMessage t;
        t <- mod_1045.get(0);
        mod_1046.put(0, t);
    endrule
    rule rule_1344;
        ChannelMessage t;
        t <- mod_1049.get(0);
        mod_1037.put(1, t);
    endrule
    rule rule_1345;
        ChannelMessage t;
        t <- mod_1041.get(1);
        mod_1042.put(1, t);
    endrule
    rule rule_1346;
        ChannelMessage t;
        t <- mod_1031.get(1);
        mod_1032.put(0, t);
    endrule
    rule rule_1347;
        ChannelMessage t;
        t <- mod_1046.get(0);
        mod_1045.put(1, t);
    endrule
    rule rule_1348;
        ChannelMessage t;
        t <- mod_1029.get(1);
        mod_1030.put(0, t);
    endrule
    rule rule_1349;
        ChannelMessage t;
        t <- mod_1032.get(1);
        mod_1033.put(0, t);
    endrule
    rule rule_1350;
        ChannelMessage t;
        t <- mod_1043.get(1);
        mod_1041.put(1, t);
    endrule
    rule rule_1351;
        ChannelMessage t;
        t <- mod_1051.get(0);
        mod_1050.put(0, t);
    endrule
    rule rule_1352;
        ChannelMessage t;
        t <- mod_1041.get(0);
        mod_1043.put(0, t);
    endrule
    rule rule_1353;
        ChannelMessage t;
        t <- mod_1034.get(0);
        mod_1035.put(0, t);
    endrule
    rule rule_1354;
        ChannelMessage t;
        t <- mod_1033.get(1);
        mod_1034.put(0, t);
    endrule
    rule rule_1355;
        ChannelMessage t;
        t <- mod_1061.get(0);
        mod_1059.put(0, t);
    endrule
    rule rule_1356;
        ChannelMessage t;
        t <- mod_1029.get(0);
        mod_1065.put(0, t);
    endrule
    rule rule_1357;
        ChannelMessage t;
        t <- mod_1026.get(0);
        mod_1027.put(0, t);
    endrule
    rule rule_1358;
        ChannelMessage t;
        t <- mod_1043.get(0);
        mod_1043.put(1, t);
    endrule
    rule rule_1359;
        ChannelMessage t;
        t <- mod_1053.get(0);
        mod_1054.put(0, t);
    endrule
    rule rule_1360;
        ChannelMessage t;
        t <- mod_1031.get(0);
        mod_1064.put(0, t);
    endrule
    rule rule_1361;
        ChannelMessage t;
        t <- mod_1040.get(1);
        mod_1041.put(0, t);
    endrule
    rule rule_1362;
        ChannelMessage t;
        t <- mod_1028.get(0);
        mod_1029.put(0, t);
    endrule
    rule rule_1363;
        ChannelMessage t;
        t <- mod_1048.get(0);
        mod_1047.put(0, t);
    endrule
    rule rule_1364;
        ChannelMessage t;
        t <- mod_1044.get(0);
        mod_1044.put(1, t);
    endrule
    rule rule_1365;
        ChannelMessage t;
        t <- mod_1055.get(0);
        mod_1053.put(0, t);
    endrule
    rule rule_1366;
        ChannelMessage t;
        t <- mod_1065.get(1);
        mod_1029.put(1, t);
    endrule
    rule rule_1367;
        ChannelMessage t;
        t <- mod_1033.get(0);
        mod_1063.put(0, t);
    endrule
    rule rule_1368;
        ChannelMessage t;
        t <- mod_1060.get(0);
        mod_1059.put(1, t);
    endrule
    rule rule_1369;
        ChannelMessage t;
        t <- mod_1036.get(0);
        mod_1037.put(0, t);
    endrule
    rule rule_1370;
        ChannelMessage t;
        t <- mod_1053.get(1);
        mod_1052.put(1, t);
    endrule
    rule rule_1371;
        ChannelMessage t;
        t <- mod_1057.get(1);
        mod_1052.put(0, t);
    endrule
    rule rule_1372;
        ChannelMessage t;
        t <- mod_1058.get(0);
        mod_1057.put(1, t);
    endrule
    rule rule_1373;
        ChannelMessage t;
        t <- mod_1027.get(0);
        mod_1028.put(0, t);
    endrule
    rule rule_1374;
        ChannelMessage t;
        t <- mod_1035.get(0);
        mod_1036.put(0, t);
    endrule
    rule rule_1375;
        ChannelMessage t;
        t <- mod_1047.get(0);
        mod_1045.put(0, t);
    endrule
    rule rule_1376;
        ChannelMessage t;
        t <- mod_1057.get(0);
        mod_1058.put(0, t);
    endrule
    rule rule_1377;
        ChannelMessage t;
        t <- mod_1063.get(0);
        mod_1033.put(1, t);
    endrule
    rule rule_1378;
        ChannelMessage t;
        t <- mod_1045.get(1);
        mod_1038.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1026.put(0, t);
        end
        if (i == 1) begin
            mod_1042.put(0, t);
        end
        if (i == 2) begin
            mod_1048.put(0, t);
        end
        if (i == 3) begin
            mod_1056.put(0, t);
        end
        if (i == 4) begin
            mod_1062.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_1030.get(0);
        end
        if (i == 3) begin
            t <- mod_1030.get(1);
        end
        if (i == 1) begin
            t <- mod_1030.get(2);
        end
        if (i == 2) begin
            t <- mod_1042.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6060 (Operation_IFC);
    Operation_IFC mod_1067_inner <- mkReshape(2, 64);
    Operation_IFC mod_1067 <- mkDebugOperation(mod_1067_inner, "mod_1067");
    Operation_IFC mod_1068_inner <- mkFlatten(1);
    Operation_IFC mod_1068 <- mkDebugOperation(mod_1068_inner, "mod_1068");
    Operation_IFC mod_1069_inner <- mkFlatten(2);
    Operation_IFC mod_1069 <- mkDebugOperation(mod_1069_inner, "mod_1069");
    Operation_IFC mod_1070_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1070 <- mkDebugOperation(mod_1070_inner, "mod_1070");
    Broadcast_IFC#(4) mod_1071_inner <- mkBroadcast(4);
    Operation_IFC mod_1071 <- mkDebugOperation(mod_1071_inner.op, "mod_1071");
    PMU_IFC mod_1072_bufferize <- mkPMU(2);
    Operation_IFC mod_1072_inner = mod_1072_bufferize.operation;
    Operation_IFC mod_1072 <- mkDebugOperation(mod_1072_inner, "mod_1072");
    Broadcast_IFC#(2) mod_1073_inner <- mkBroadcast(2);
    Operation_IFC mod_1073 <- mkDebugOperation(mod_1073_inner.op, "mod_1073");
    PMU_IFC mod_1074_bufferize <- mkPMU(1);
    Operation_IFC mod_1074_inner = mod_1074_bufferize.operation;
    Operation_IFC mod_1074 <- mkDebugOperation(mod_1074_inner, "mod_1074");
    Operation_IFC mod_1075_inner <- mkBinaryMap(1130, matmul_t_tile);
    Operation_IFC mod_1075 <- mkDebugOperation(mod_1075_inner, "mod_1075");
    Operation_IFC mod_1076_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1076 <- mkDebugOperation(mod_1076_inner, "mod_1076");
    Operation_IFC mod_1077_inner <- mkBinaryMap(1898, mul_tile);
    Operation_IFC mod_1077 <- mkDebugOperation(mod_1077_inner, "mod_1077");
    PMU_IFC mod_1078_bufferize <- mkPMU(1);
    Operation_IFC mod_1078_inner = mod_1078_bufferize.operation;
    Operation_IFC mod_1078 <- mkDebugOperation(mod_1078_inner, "mod_1078");
    Operation_IFC mod_1079_inner <- mkBinaryMap(2511, matmul_t_tile);
    Operation_IFC mod_1079 <- mkDebugOperation(mod_1079_inner, "mod_1079");
    Operation_IFC mod_1080_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1080 <- mkDebugOperation(mod_1080_inner, "mod_1080");
    Operation_IFC mod_1081_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1081 <- mkDebugOperation(mod_1081_inner, "mod_1081");
    Operation_IFC mod_1082_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1082 <- mkDebugOperation(mod_1082_inner, "mod_1082");
    Operation_IFC mod_1083_inner <- mkBinaryMap(2797, mul_tile);
    Operation_IFC mod_1083 <- mkDebugOperation(mod_1083_inner, "mod_1083");
    PMU_IFC mod_1084_bufferize <- mkPMU(1);
    Operation_IFC mod_1084_inner = mod_1084_bufferize.operation;
    Operation_IFC mod_1084 <- mkDebugOperation(mod_1084_inner, "mod_1084");
    PMU_IFC mod_1085_bufferize <- mkPMU(2);
    Operation_IFC mod_1085_inner = mod_1085_bufferize.operation;
    Operation_IFC mod_1085 <- mkDebugOperation(mod_1085_inner, "mod_1085");
    PMU_IFC mod_1086_bufferize <- mkPMU(2);
    Operation_IFC mod_1086_inner = mod_1086_bufferize.operation;
    Operation_IFC mod_1086 <- mkDebugOperation(mod_1086_inner, "mod_1086");
    Operation_IFC mod_1087_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1087 <- mkDebugOperation(mod_1087_inner, "mod_1087");
    Operation_IFC mod_1088_inner <- mkFlatten(1);
    Operation_IFC mod_1088 <- mkDebugOperation(mod_1088_inner, "mod_1088");
    Operation_IFC mod_1089_inner <- mkFlatten(0);
    Operation_IFC mod_1089 <- mkDebugOperation(mod_1089_inner, "mod_1089");
    Operation_IFC mod_1090_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1090 <- mkDebugOperation(mod_1090_inner, "mod_1090");
    Operation_IFC mod_1091_inner <- mkUnaryMap(1770, silu_tile);
    Operation_IFC mod_1091 <- mkDebugOperation(mod_1091_inner, "mod_1091");
    Operation_IFC mod_1092_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1092 <- mkDebugOperation(mod_1092_inner, "mod_1092");
    Operation_IFC mod_1093_inner <- mkBinaryMap(1642, matmul_t_tile);
    Operation_IFC mod_1093 <- mkDebugOperation(mod_1093_inner, "mod_1093");
    PMU_IFC mod_1094_bufferize <- mkPMU(2);
    Operation_IFC mod_1094_inner = mod_1094_bufferize.operation;
    Operation_IFC mod_1094 <- mkDebugOperation(mod_1094_inner, "mod_1094");
    Operation_IFC mod_1095_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1095 <- mkDebugOperation(mod_1095_inner, "mod_1095");
    Operation_IFC mod_1096_inner <- mkFlatten(1);
    Operation_IFC mod_1096 <- mkDebugOperation(mod_1096_inner, "mod_1096");
    Operation_IFC mod_1097_inner <- mkFlatten(0);
    Operation_IFC mod_1097 <- mkDebugOperation(mod_1097_inner, "mod_1097");
    PMU_IFC mod_1098_bufferize <- mkPMU(1);
    Operation_IFC mod_1098_inner = mod_1098_bufferize.operation;
    Operation_IFC mod_1098 <- mkDebugOperation(mod_1098_inner, "mod_1098");
    Operation_IFC mod_1099_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1099 <- mkDebugOperation(mod_1099_inner, "mod_1099");
    PMU_IFC mod_1100_bufferize <- mkPMU(2);
    Operation_IFC mod_1100_inner = mod_1100_bufferize.operation;
    Operation_IFC mod_1100 <- mkDebugOperation(mod_1100_inner, "mod_1100");
    Operation_IFC mod_1101_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1101 <- mkDebugOperation(mod_1101_inner, "mod_1101");
    Operation_IFC mod_1102_inner <- mkFlatten(1);
    Operation_IFC mod_1102 <- mkDebugOperation(mod_1102_inner, "mod_1102");
    Operation_IFC mod_1103_inner <- mkFlatten(0);
    Operation_IFC mod_1103 <- mkDebugOperation(mod_1103_inner, "mod_1103");
    Operation_IFC mod_1104_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1104 <- mkDebugOperation(mod_1104_inner, "mod_1104");
    Operation_IFC mod_1105_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1105 <- mkDebugOperation(mod_1105_inner, "mod_1105");
    PMU_IFC mod_1106_bufferize <- mkPMU(2);
    Operation_IFC mod_1106_inner = mod_1106_bufferize.operation;
    Operation_IFC mod_1106 <- mkDebugOperation(mod_1106_inner, "mod_1106");
    rule rule_1379;
        ChannelMessage t;
        t <- mod_1078.get(0);
        mod_1090.put(0, t);
    endrule
    rule rule_1380;
        ChannelMessage t;
        t <- mod_1085.get(0);
        mod_1085.put(1, t);
    endrule
    rule rule_1381;
        ChannelMessage t;
        t <- mod_1077.get(0);
        mod_1078.put(0, t);
    endrule
    rule rule_1382;
        ChannelMessage t;
        t <- mod_1086.get(1);
        mod_1079.put(1, t);
    endrule
    rule rule_1383;
        ChannelMessage t;
        t <- mod_1084.get(0);
        mod_1084.put(1, t);
    endrule
    rule rule_1384;
        ChannelMessage t;
        t <- mod_1090.get(0);
        mod_1078.put(1, t);
    endrule
    rule rule_1385;
        ChannelMessage t;
        t <- mod_1092.get(0);
        mod_1091.put(0, t);
    endrule
    rule rule_1386;
        ChannelMessage t;
        t <- mod_1074.get(1);
        mod_1075.put(0, t);
    endrule
    rule rule_1387;
        ChannelMessage t;
        t <- mod_1069.get(0);
        mod_1070.put(0, t);
    endrule
    rule rule_1388;
        ChannelMessage t;
        t <- mod_1080.get(0);
        mod_1081.put(0, t);
    endrule
    rule rule_1389;
        ChannelMessage t;
        t <- mod_1079.get(0);
        mod_1080.put(0, t);
    endrule
    rule rule_1390;
        ChannelMessage t;
        t <- mod_1076.get(0);
        mod_1077.put(0, t);
    endrule
    rule rule_1391;
        ChannelMessage t;
        t <- mod_1071.get(3);
        mod_1072.put(0, t);
    endrule
    rule rule_1392;
        ChannelMessage t;
        t <- mod_1091.get(0);
        mod_1077.put(1, t);
    endrule
    rule rule_1393;
        ChannelMessage t;
        t <- mod_1097.get(0);
        mod_1096.put(0, t);
    endrule
    rule rule_1394;
        ChannelMessage t;
        t <- mod_1072.get(1);
        mod_1073.put(0, t);
    endrule
    rule rule_1395;
        ChannelMessage t;
        t <- mod_1094.get(1);
        mod_1093.put(1, t);
    endrule
    rule rule_1396;
        ChannelMessage t;
        t <- mod_1098.get(0);
        mod_1099.put(0, t);
    endrule
    rule rule_1397;
        ChannelMessage t;
        t <- mod_1104.get(0);
        mod_1074.put(1, t);
    endrule
    rule rule_1398;
        ChannelMessage t;
        t <- mod_1070.get(1);
        mod_1071.put(0, t);
    endrule
    rule rule_1399;
        ChannelMessage t;
        t <- mod_1067.get(0);
        mod_1068.put(0, t);
    endrule
    rule rule_1400;
        ChannelMessage t;
        t <- mod_1073.get(1);
        mod_1074.put(0, t);
    endrule
    rule rule_1401;
        ChannelMessage t;
        t <- mod_1096.get(0);
        mod_1094.put(0, t);
    endrule
    rule rule_1402;
        ChannelMessage t;
        t <- mod_1084.get(1);
        mod_1082.put(1, t);
    endrule
    rule rule_1403;
        ChannelMessage t;
        t <- mod_1098.get(1);
        mod_1093.put(0, t);
    endrule
    rule rule_1404;
        ChannelMessage t;
        t <- mod_1081.get(1);
        mod_1082.put(0, t);
    endrule
    rule rule_1405;
        ChannelMessage t;
        t <- mod_1074.get(0);
        mod_1104.put(0, t);
    endrule
    rule rule_1406;
        ChannelMessage t;
        t <- mod_1082.get(0);
        mod_1084.put(0, t);
    endrule
    rule rule_1407;
        ChannelMessage t;
        t <- mod_1101.get(0);
        mod_1100.put(1, t);
    endrule
    rule rule_1408;
        ChannelMessage t;
        t <- mod_1088.get(0);
        mod_1086.put(0, t);
    endrule
    rule rule_1409;
        ChannelMessage t;
        t <- mod_1103.get(0);
        mod_1102.put(0, t);
    endrule
    rule rule_1410;
        ChannelMessage t;
        t <- mod_1106.get(0);
        mod_1106.put(1, t);
    endrule
    rule rule_1411;
        ChannelMessage t;
        t <- mod_1106.get(1);
        mod_1070.put(1, t);
    endrule
    rule rule_1412;
        ChannelMessage t;
        t <- mod_1099.get(0);
        mod_1098.put(1, t);
    endrule
    rule rule_1413;
        ChannelMessage t;
        t <- mod_1081.get(0);
        mod_1085.put(0, t);
    endrule
    rule rule_1414;
        ChannelMessage t;
        t <- mod_1089.get(0);
        mod_1088.put(0, t);
    endrule
    rule rule_1415;
        ChannelMessage t;
        t <- mod_1087.get(0);
        mod_1086.put(1, t);
    endrule
    rule rule_1416;
        ChannelMessage t;
        t <- mod_1072.get(0);
        mod_1105.put(0, t);
    endrule
    rule rule_1417;
        ChannelMessage t;
        t <- mod_1100.get(1);
        mod_1075.put(1, t);
    endrule
    rule rule_1418;
        ChannelMessage t;
        t <- mod_1073.get(0);
        mod_1098.put(0, t);
    endrule
    rule rule_1419;
        ChannelMessage t;
        t <- mod_1100.get(0);
        mod_1101.put(0, t);
    endrule
    rule rule_1420;
        ChannelMessage t;
        t <- mod_1085.get(1);
        mod_1081.put(1, t);
    endrule
    rule rule_1421;
        ChannelMessage t;
        t <- mod_1078.get(1);
        mod_1079.put(0, t);
    endrule
    rule rule_1422;
        ChannelMessage t;
        t <- mod_1105.get(0);
        mod_1072.put(1, t);
    endrule
    rule rule_1423;
        ChannelMessage t;
        t <- mod_1095.get(0);
        mod_1094.put(1, t);
    endrule
    rule rule_1424;
        ChannelMessage t;
        t <- mod_1094.get(0);
        mod_1095.put(0, t);
    endrule
    rule rule_1425;
        ChannelMessage t;
        t <- mod_1086.get(0);
        mod_1087.put(0, t);
    endrule
    rule rule_1426;
        ChannelMessage t;
        t <- mod_1102.get(0);
        mod_1100.put(0, t);
    endrule
    rule rule_1427;
        ChannelMessage t;
        t <- mod_1075.get(0);
        mod_1076.put(0, t);
    endrule
    rule rule_1428;
        ChannelMessage t;
        t <- mod_1093.get(0);
        mod_1092.put(0, t);
    endrule
    rule rule_1429;
        ChannelMessage t;
        t <- mod_1082.get(1);
        mod_1083.put(1, t);
    endrule
    rule rule_1430;
        ChannelMessage t;
        t <- mod_1068.get(0);
        mod_1069.put(0, t);
    endrule
    rule rule_1431;
        ChannelMessage t;
        t <- mod_1070.get(0);
        mod_1106.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1067.put(0, t);
        end
        if (i == 1) begin
            mod_1083.put(0, t);
        end
        if (i == 2) begin
            mod_1089.put(0, t);
        end
        if (i == 3) begin
            mod_1097.put(0, t);
        end
        if (i == 4) begin
            mod_1103.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_1071.get(0);
        end
        if (i == 0) begin
            t <- mod_1071.get(1);
        end
        if (i == 2) begin
            t <- mod_1071.get(2);
        end
        if (i == 1) begin
            t <- mod_1083.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6061 (Operation_IFC);
    Operation_IFC mod_1108_inner <- mkReshape(2, 64);
    Operation_IFC mod_1108 <- mkDebugOperation(mod_1108_inner, "mod_1108");
    Operation_IFC mod_1109_inner <- mkFlatten(1);
    Operation_IFC mod_1109 <- mkDebugOperation(mod_1109_inner, "mod_1109");
    Operation_IFC mod_1110_inner <- mkFlatten(2);
    Operation_IFC mod_1110 <- mkDebugOperation(mod_1110_inner, "mod_1110");
    Operation_IFC mod_1111_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1111 <- mkDebugOperation(mod_1111_inner, "mod_1111");
    Broadcast_IFC#(4) mod_1112_inner <- mkBroadcast(4);
    Operation_IFC mod_1112 <- mkDebugOperation(mod_1112_inner.op, "mod_1112");
    PMU_IFC mod_1113_bufferize <- mkPMU(2);
    Operation_IFC mod_1113_inner = mod_1113_bufferize.operation;
    Operation_IFC mod_1113 <- mkDebugOperation(mod_1113_inner, "mod_1113");
    Broadcast_IFC#(2) mod_1114_inner <- mkBroadcast(2);
    Operation_IFC mod_1114 <- mkDebugOperation(mod_1114_inner.op, "mod_1114");
    PMU_IFC mod_1115_bufferize <- mkPMU(1);
    Operation_IFC mod_1115_inner = mod_1115_bufferize.operation;
    Operation_IFC mod_1115 <- mkDebugOperation(mod_1115_inner, "mod_1115");
    Operation_IFC mod_1116_inner <- mkBinaryMap(1129, matmul_t_tile);
    Operation_IFC mod_1116 <- mkDebugOperation(mod_1116_inner, "mod_1116");
    Operation_IFC mod_1117_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1117 <- mkDebugOperation(mod_1117_inner, "mod_1117");
    Operation_IFC mod_1118_inner <- mkBinaryMap(1897, mul_tile);
    Operation_IFC mod_1118 <- mkDebugOperation(mod_1118_inner, "mod_1118");
    PMU_IFC mod_1119_bufferize <- mkPMU(1);
    Operation_IFC mod_1119_inner = mod_1119_bufferize.operation;
    Operation_IFC mod_1119 <- mkDebugOperation(mod_1119_inner, "mod_1119");
    Operation_IFC mod_1120_inner <- mkBinaryMap(2509, matmul_t_tile);
    Operation_IFC mod_1120 <- mkDebugOperation(mod_1120_inner, "mod_1120");
    Operation_IFC mod_1121_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1121 <- mkDebugOperation(mod_1121_inner, "mod_1121");
    Operation_IFC mod_1122_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1122 <- mkDebugOperation(mod_1122_inner, "mod_1122");
    Operation_IFC mod_1123_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1123 <- mkDebugOperation(mod_1123_inner, "mod_1123");
    Operation_IFC mod_1124_inner <- mkBinaryMap(2796, mul_tile);
    Operation_IFC mod_1124 <- mkDebugOperation(mod_1124_inner, "mod_1124");
    PMU_IFC mod_1125_bufferize <- mkPMU(1);
    Operation_IFC mod_1125_inner = mod_1125_bufferize.operation;
    Operation_IFC mod_1125 <- mkDebugOperation(mod_1125_inner, "mod_1125");
    PMU_IFC mod_1126_bufferize <- mkPMU(2);
    Operation_IFC mod_1126_inner = mod_1126_bufferize.operation;
    Operation_IFC mod_1126 <- mkDebugOperation(mod_1126_inner, "mod_1126");
    PMU_IFC mod_1127_bufferize <- mkPMU(2);
    Operation_IFC mod_1127_inner = mod_1127_bufferize.operation;
    Operation_IFC mod_1127 <- mkDebugOperation(mod_1127_inner, "mod_1127");
    Operation_IFC mod_1128_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1128 <- mkDebugOperation(mod_1128_inner, "mod_1128");
    Operation_IFC mod_1129_inner <- mkFlatten(1);
    Operation_IFC mod_1129 <- mkDebugOperation(mod_1129_inner, "mod_1129");
    Operation_IFC mod_1130_inner <- mkFlatten(0);
    Operation_IFC mod_1130 <- mkDebugOperation(mod_1130_inner, "mod_1130");
    Operation_IFC mod_1131_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1131 <- mkDebugOperation(mod_1131_inner, "mod_1131");
    Operation_IFC mod_1132_inner <- mkUnaryMap(1769, silu_tile);
    Operation_IFC mod_1132 <- mkDebugOperation(mod_1132_inner, "mod_1132");
    Operation_IFC mod_1133_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1133 <- mkDebugOperation(mod_1133_inner, "mod_1133");
    Operation_IFC mod_1134_inner <- mkBinaryMap(1641, matmul_t_tile);
    Operation_IFC mod_1134 <- mkDebugOperation(mod_1134_inner, "mod_1134");
    PMU_IFC mod_1135_bufferize <- mkPMU(2);
    Operation_IFC mod_1135_inner = mod_1135_bufferize.operation;
    Operation_IFC mod_1135 <- mkDebugOperation(mod_1135_inner, "mod_1135");
    Operation_IFC mod_1136_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1136 <- mkDebugOperation(mod_1136_inner, "mod_1136");
    Operation_IFC mod_1137_inner <- mkFlatten(1);
    Operation_IFC mod_1137 <- mkDebugOperation(mod_1137_inner, "mod_1137");
    Operation_IFC mod_1138_inner <- mkFlatten(0);
    Operation_IFC mod_1138 <- mkDebugOperation(mod_1138_inner, "mod_1138");
    PMU_IFC mod_1139_bufferize <- mkPMU(1);
    Operation_IFC mod_1139_inner = mod_1139_bufferize.operation;
    Operation_IFC mod_1139 <- mkDebugOperation(mod_1139_inner, "mod_1139");
    Operation_IFC mod_1140_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1140 <- mkDebugOperation(mod_1140_inner, "mod_1140");
    PMU_IFC mod_1141_bufferize <- mkPMU(2);
    Operation_IFC mod_1141_inner = mod_1141_bufferize.operation;
    Operation_IFC mod_1141 <- mkDebugOperation(mod_1141_inner, "mod_1141");
    Operation_IFC mod_1142_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1142 <- mkDebugOperation(mod_1142_inner, "mod_1142");
    Operation_IFC mod_1143_inner <- mkFlatten(1);
    Operation_IFC mod_1143 <- mkDebugOperation(mod_1143_inner, "mod_1143");
    Operation_IFC mod_1144_inner <- mkFlatten(0);
    Operation_IFC mod_1144 <- mkDebugOperation(mod_1144_inner, "mod_1144");
    Operation_IFC mod_1145_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1145 <- mkDebugOperation(mod_1145_inner, "mod_1145");
    Operation_IFC mod_1146_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1146 <- mkDebugOperation(mod_1146_inner, "mod_1146");
    PMU_IFC mod_1147_bufferize <- mkPMU(2);
    Operation_IFC mod_1147_inner = mod_1147_bufferize.operation;
    Operation_IFC mod_1147 <- mkDebugOperation(mod_1147_inner, "mod_1147");
    rule rule_1432;
        ChannelMessage t;
        t <- mod_1135.get(0);
        mod_1136.put(0, t);
    endrule
    rule rule_1433;
        ChannelMessage t;
        t <- mod_1134.get(0);
        mod_1133.put(0, t);
    endrule
    rule rule_1434;
        ChannelMessage t;
        t <- mod_1117.get(0);
        mod_1118.put(0, t);
    endrule
    rule rule_1435;
        ChannelMessage t;
        t <- mod_1136.get(0);
        mod_1135.put(1, t);
    endrule
    rule rule_1436;
        ChannelMessage t;
        t <- mod_1130.get(0);
        mod_1129.put(0, t);
    endrule
    rule rule_1437;
        ChannelMessage t;
        t <- mod_1141.get(0);
        mod_1142.put(0, t);
    endrule
    rule rule_1438;
        ChannelMessage t;
        t <- mod_1142.get(0);
        mod_1141.put(1, t);
    endrule
    rule rule_1439;
        ChannelMessage t;
        t <- mod_1113.get(1);
        mod_1114.put(0, t);
    endrule
    rule rule_1440;
        ChannelMessage t;
        t <- mod_1115.get(1);
        mod_1116.put(0, t);
    endrule
    rule rule_1441;
        ChannelMessage t;
        t <- mod_1147.get(0);
        mod_1147.put(1, t);
    endrule
    rule rule_1442;
        ChannelMessage t;
        t <- mod_1127.get(0);
        mod_1128.put(0, t);
    endrule
    rule rule_1443;
        ChannelMessage t;
        t <- mod_1120.get(0);
        mod_1121.put(0, t);
    endrule
    rule rule_1444;
        ChannelMessage t;
        t <- mod_1123.get(1);
        mod_1124.put(1, t);
    endrule
    rule rule_1445;
        ChannelMessage t;
        t <- mod_1141.get(1);
        mod_1116.put(1, t);
    endrule
    rule rule_1446;
        ChannelMessage t;
        t <- mod_1131.get(0);
        mod_1119.put(1, t);
    endrule
    rule rule_1447;
        ChannelMessage t;
        t <- mod_1143.get(0);
        mod_1141.put(0, t);
    endrule
    rule rule_1448;
        ChannelMessage t;
        t <- mod_1127.get(1);
        mod_1120.put(1, t);
    endrule
    rule rule_1449;
        ChannelMessage t;
        t <- mod_1133.get(0);
        mod_1132.put(0, t);
    endrule
    rule rule_1450;
        ChannelMessage t;
        t <- mod_1125.get(1);
        mod_1123.put(1, t);
    endrule
    rule rule_1451;
        ChannelMessage t;
        t <- mod_1108.get(0);
        mod_1109.put(0, t);
    endrule
    rule rule_1452;
        ChannelMessage t;
        t <- mod_1118.get(0);
        mod_1119.put(0, t);
    endrule
    rule rule_1453;
        ChannelMessage t;
        t <- mod_1119.get(1);
        mod_1120.put(0, t);
    endrule
    rule rule_1454;
        ChannelMessage t;
        t <- mod_1110.get(0);
        mod_1111.put(0, t);
    endrule
    rule rule_1455;
        ChannelMessage t;
        t <- mod_1140.get(0);
        mod_1139.put(1, t);
    endrule
    rule rule_1456;
        ChannelMessage t;
        t <- mod_1147.get(1);
        mod_1111.put(1, t);
    endrule
    rule rule_1457;
        ChannelMessage t;
        t <- mod_1123.get(0);
        mod_1125.put(0, t);
    endrule
    rule rule_1458;
        ChannelMessage t;
        t <- mod_1114.get(1);
        mod_1115.put(0, t);
    endrule
    rule rule_1459;
        ChannelMessage t;
        t <- mod_1109.get(0);
        mod_1110.put(0, t);
    endrule
    rule rule_1460;
        ChannelMessage t;
        t <- mod_1126.get(0);
        mod_1126.put(1, t);
    endrule
    rule rule_1461;
        ChannelMessage t;
        t <- mod_1111.get(1);
        mod_1112.put(0, t);
    endrule
    rule rule_1462;
        ChannelMessage t;
        t <- mod_1125.get(0);
        mod_1125.put(1, t);
    endrule
    rule rule_1463;
        ChannelMessage t;
        t <- mod_1144.get(0);
        mod_1143.put(0, t);
    endrule
    rule rule_1464;
        ChannelMessage t;
        t <- mod_1122.get(1);
        mod_1123.put(0, t);
    endrule
    rule rule_1465;
        ChannelMessage t;
        t <- mod_1146.get(0);
        mod_1113.put(1, t);
    endrule
    rule rule_1466;
        ChannelMessage t;
        t <- mod_1137.get(0);
        mod_1135.put(0, t);
    endrule
    rule rule_1467;
        ChannelMessage t;
        t <- mod_1132.get(0);
        mod_1118.put(1, t);
    endrule
    rule rule_1468;
        ChannelMessage t;
        t <- mod_1114.get(0);
        mod_1139.put(0, t);
    endrule
    rule rule_1469;
        ChannelMessage t;
        t <- mod_1139.get(0);
        mod_1140.put(0, t);
    endrule
    rule rule_1470;
        ChannelMessage t;
        t <- mod_1128.get(0);
        mod_1127.put(1, t);
    endrule
    rule rule_1471;
        ChannelMessage t;
        t <- mod_1126.get(1);
        mod_1122.put(1, t);
    endrule
    rule rule_1472;
        ChannelMessage t;
        t <- mod_1111.get(0);
        mod_1147.put(0, t);
    endrule
    rule rule_1473;
        ChannelMessage t;
        t <- mod_1112.get(3);
        mod_1113.put(0, t);
    endrule
    rule rule_1474;
        ChannelMessage t;
        t <- mod_1115.get(0);
        mod_1145.put(0, t);
    endrule
    rule rule_1475;
        ChannelMessage t;
        t <- mod_1122.get(0);
        mod_1126.put(0, t);
    endrule
    rule rule_1476;
        ChannelMessage t;
        t <- mod_1145.get(0);
        mod_1115.put(1, t);
    endrule
    rule rule_1477;
        ChannelMessage t;
        t <- mod_1119.get(0);
        mod_1131.put(0, t);
    endrule
    rule rule_1478;
        ChannelMessage t;
        t <- mod_1135.get(1);
        mod_1134.put(1, t);
    endrule
    rule rule_1479;
        ChannelMessage t;
        t <- mod_1138.get(0);
        mod_1137.put(0, t);
    endrule
    rule rule_1480;
        ChannelMessage t;
        t <- mod_1139.get(1);
        mod_1134.put(0, t);
    endrule
    rule rule_1481;
        ChannelMessage t;
        t <- mod_1129.get(0);
        mod_1127.put(0, t);
    endrule
    rule rule_1482;
        ChannelMessage t;
        t <- mod_1113.get(0);
        mod_1146.put(0, t);
    endrule
    rule rule_1483;
        ChannelMessage t;
        t <- mod_1121.get(0);
        mod_1122.put(0, t);
    endrule
    rule rule_1484;
        ChannelMessage t;
        t <- mod_1116.get(0);
        mod_1117.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1108.put(0, t);
        end
        if (i == 1) begin
            mod_1124.put(0, t);
        end
        if (i == 2) begin
            mod_1130.put(0, t);
        end
        if (i == 3) begin
            mod_1138.put(0, t);
        end
        if (i == 4) begin
            mod_1144.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_1112.get(0);
        end
        if (i == 0) begin
            t <- mod_1112.get(1);
        end
        if (i == 3) begin
            t <- mod_1112.get(2);
        end
        if (i == 2) begin
            t <- mod_1124.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6062 (Operation_IFC);
    Operation_IFC mod_1149_inner <- mkReshape(2, 64);
    Operation_IFC mod_1149 <- mkDebugOperation(mod_1149_inner, "mod_1149");
    Operation_IFC mod_1150_inner <- mkFlatten(1);
    Operation_IFC mod_1150 <- mkDebugOperation(mod_1150_inner, "mod_1150");
    Operation_IFC mod_1151_inner <- mkFlatten(2);
    Operation_IFC mod_1151 <- mkDebugOperation(mod_1151_inner, "mod_1151");
    Operation_IFC mod_1152_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1152 <- mkDebugOperation(mod_1152_inner, "mod_1152");
    Broadcast_IFC#(4) mod_1153_inner <- mkBroadcast(4);
    Operation_IFC mod_1153 <- mkDebugOperation(mod_1153_inner.op, "mod_1153");
    PMU_IFC mod_1154_bufferize <- mkPMU(2);
    Operation_IFC mod_1154_inner = mod_1154_bufferize.operation;
    Operation_IFC mod_1154 <- mkDebugOperation(mod_1154_inner, "mod_1154");
    Broadcast_IFC#(2) mod_1155_inner <- mkBroadcast(2);
    Operation_IFC mod_1155 <- mkDebugOperation(mod_1155_inner.op, "mod_1155");
    PMU_IFC mod_1156_bufferize <- mkPMU(1);
    Operation_IFC mod_1156_inner = mod_1156_bufferize.operation;
    Operation_IFC mod_1156 <- mkDebugOperation(mod_1156_inner, "mod_1156");
    Operation_IFC mod_1157_inner <- mkBinaryMap(1128, matmul_t_tile);
    Operation_IFC mod_1157 <- mkDebugOperation(mod_1157_inner, "mod_1157");
    Operation_IFC mod_1158_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1158 <- mkDebugOperation(mod_1158_inner, "mod_1158");
    Operation_IFC mod_1159_inner <- mkBinaryMap(1896, mul_tile);
    Operation_IFC mod_1159 <- mkDebugOperation(mod_1159_inner, "mod_1159");
    PMU_IFC mod_1160_bufferize <- mkPMU(1);
    Operation_IFC mod_1160_inner = mod_1160_bufferize.operation;
    Operation_IFC mod_1160 <- mkDebugOperation(mod_1160_inner, "mod_1160");
    Operation_IFC mod_1161_inner <- mkBinaryMap(2507, matmul_t_tile);
    Operation_IFC mod_1161 <- mkDebugOperation(mod_1161_inner, "mod_1161");
    Operation_IFC mod_1162_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1162 <- mkDebugOperation(mod_1162_inner, "mod_1162");
    Operation_IFC mod_1163_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1163 <- mkDebugOperation(mod_1163_inner, "mod_1163");
    Operation_IFC mod_1164_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1164 <- mkDebugOperation(mod_1164_inner, "mod_1164");
    Operation_IFC mod_1165_inner <- mkBinaryMap(2795, mul_tile);
    Operation_IFC mod_1165 <- mkDebugOperation(mod_1165_inner, "mod_1165");
    PMU_IFC mod_1166_bufferize <- mkPMU(1);
    Operation_IFC mod_1166_inner = mod_1166_bufferize.operation;
    Operation_IFC mod_1166 <- mkDebugOperation(mod_1166_inner, "mod_1166");
    PMU_IFC mod_1167_bufferize <- mkPMU(2);
    Operation_IFC mod_1167_inner = mod_1167_bufferize.operation;
    Operation_IFC mod_1167 <- mkDebugOperation(mod_1167_inner, "mod_1167");
    PMU_IFC mod_1168_bufferize <- mkPMU(2);
    Operation_IFC mod_1168_inner = mod_1168_bufferize.operation;
    Operation_IFC mod_1168 <- mkDebugOperation(mod_1168_inner, "mod_1168");
    Operation_IFC mod_1169_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1169 <- mkDebugOperation(mod_1169_inner, "mod_1169");
    Operation_IFC mod_1170_inner <- mkFlatten(1);
    Operation_IFC mod_1170 <- mkDebugOperation(mod_1170_inner, "mod_1170");
    Operation_IFC mod_1171_inner <- mkFlatten(0);
    Operation_IFC mod_1171 <- mkDebugOperation(mod_1171_inner, "mod_1171");
    Operation_IFC mod_1172_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1172 <- mkDebugOperation(mod_1172_inner, "mod_1172");
    Operation_IFC mod_1173_inner <- mkUnaryMap(1768, silu_tile);
    Operation_IFC mod_1173 <- mkDebugOperation(mod_1173_inner, "mod_1173");
    Operation_IFC mod_1174_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1174 <- mkDebugOperation(mod_1174_inner, "mod_1174");
    Operation_IFC mod_1175_inner <- mkBinaryMap(1640, matmul_t_tile);
    Operation_IFC mod_1175 <- mkDebugOperation(mod_1175_inner, "mod_1175");
    PMU_IFC mod_1176_bufferize <- mkPMU(2);
    Operation_IFC mod_1176_inner = mod_1176_bufferize.operation;
    Operation_IFC mod_1176 <- mkDebugOperation(mod_1176_inner, "mod_1176");
    Operation_IFC mod_1177_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1177 <- mkDebugOperation(mod_1177_inner, "mod_1177");
    Operation_IFC mod_1178_inner <- mkFlatten(1);
    Operation_IFC mod_1178 <- mkDebugOperation(mod_1178_inner, "mod_1178");
    Operation_IFC mod_1179_inner <- mkFlatten(0);
    Operation_IFC mod_1179 <- mkDebugOperation(mod_1179_inner, "mod_1179");
    PMU_IFC mod_1180_bufferize <- mkPMU(1);
    Operation_IFC mod_1180_inner = mod_1180_bufferize.operation;
    Operation_IFC mod_1180 <- mkDebugOperation(mod_1180_inner, "mod_1180");
    Operation_IFC mod_1181_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1181 <- mkDebugOperation(mod_1181_inner, "mod_1181");
    PMU_IFC mod_1182_bufferize <- mkPMU(2);
    Operation_IFC mod_1182_inner = mod_1182_bufferize.operation;
    Operation_IFC mod_1182 <- mkDebugOperation(mod_1182_inner, "mod_1182");
    Operation_IFC mod_1183_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1183 <- mkDebugOperation(mod_1183_inner, "mod_1183");
    Operation_IFC mod_1184_inner <- mkFlatten(1);
    Operation_IFC mod_1184 <- mkDebugOperation(mod_1184_inner, "mod_1184");
    Operation_IFC mod_1185_inner <- mkFlatten(0);
    Operation_IFC mod_1185 <- mkDebugOperation(mod_1185_inner, "mod_1185");
    Operation_IFC mod_1186_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1186 <- mkDebugOperation(mod_1186_inner, "mod_1186");
    Operation_IFC mod_1187_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1187 <- mkDebugOperation(mod_1187_inner, "mod_1187");
    PMU_IFC mod_1188_bufferize <- mkPMU(2);
    Operation_IFC mod_1188_inner = mod_1188_bufferize.operation;
    Operation_IFC mod_1188 <- mkDebugOperation(mod_1188_inner, "mod_1188");
    rule rule_1485;
        ChannelMessage t;
        t <- mod_1160.get(0);
        mod_1172.put(0, t);
    endrule
    rule rule_1486;
        ChannelMessage t;
        t <- mod_1168.get(0);
        mod_1169.put(0, t);
    endrule
    rule rule_1487;
        ChannelMessage t;
        t <- mod_1170.get(0);
        mod_1168.put(0, t);
    endrule
    rule rule_1488;
        ChannelMessage t;
        t <- mod_1182.get(0);
        mod_1183.put(0, t);
    endrule
    rule rule_1489;
        ChannelMessage t;
        t <- mod_1156.get(1);
        mod_1157.put(0, t);
    endrule
    rule rule_1490;
        ChannelMessage t;
        t <- mod_1164.get(0);
        mod_1166.put(0, t);
    endrule
    rule rule_1491;
        ChannelMessage t;
        t <- mod_1186.get(0);
        mod_1156.put(1, t);
    endrule
    rule rule_1492;
        ChannelMessage t;
        t <- mod_1188.get(0);
        mod_1188.put(1, t);
    endrule
    rule rule_1493;
        ChannelMessage t;
        t <- mod_1152.get(0);
        mod_1188.put(0, t);
    endrule
    rule rule_1494;
        ChannelMessage t;
        t <- mod_1177.get(0);
        mod_1176.put(1, t);
    endrule
    rule rule_1495;
        ChannelMessage t;
        t <- mod_1166.get(0);
        mod_1166.put(1, t);
    endrule
    rule rule_1496;
        ChannelMessage t;
        t <- mod_1163.get(0);
        mod_1167.put(0, t);
    endrule
    rule rule_1497;
        ChannelMessage t;
        t <- mod_1180.get(0);
        mod_1181.put(0, t);
    endrule
    rule rule_1498;
        ChannelMessage t;
        t <- mod_1180.get(1);
        mod_1175.put(0, t);
    endrule
    rule rule_1499;
        ChannelMessage t;
        t <- mod_1149.get(0);
        mod_1150.put(0, t);
    endrule
    rule rule_1500;
        ChannelMessage t;
        t <- mod_1167.get(1);
        mod_1163.put(1, t);
    endrule
    rule rule_1501;
        ChannelMessage t;
        t <- mod_1156.get(0);
        mod_1186.put(0, t);
    endrule
    rule rule_1502;
        ChannelMessage t;
        t <- mod_1158.get(0);
        mod_1159.put(0, t);
    endrule
    rule rule_1503;
        ChannelMessage t;
        t <- mod_1159.get(0);
        mod_1160.put(0, t);
    endrule
    rule rule_1504;
        ChannelMessage t;
        t <- mod_1176.get(0);
        mod_1177.put(0, t);
    endrule
    rule rule_1505;
        ChannelMessage t;
        t <- mod_1155.get(1);
        mod_1156.put(0, t);
    endrule
    rule rule_1506;
        ChannelMessage t;
        t <- mod_1150.get(0);
        mod_1151.put(0, t);
    endrule
    rule rule_1507;
        ChannelMessage t;
        t <- mod_1162.get(0);
        mod_1163.put(0, t);
    endrule
    rule rule_1508;
        ChannelMessage t;
        t <- mod_1176.get(1);
        mod_1175.put(1, t);
    endrule
    rule rule_1509;
        ChannelMessage t;
        t <- mod_1166.get(1);
        mod_1164.put(1, t);
    endrule
    rule rule_1510;
        ChannelMessage t;
        t <- mod_1181.get(0);
        mod_1180.put(1, t);
    endrule
    rule rule_1511;
        ChannelMessage t;
        t <- mod_1167.get(0);
        mod_1167.put(1, t);
    endrule
    rule rule_1512;
        ChannelMessage t;
        t <- mod_1169.get(0);
        mod_1168.put(1, t);
    endrule
    rule rule_1513;
        ChannelMessage t;
        t <- mod_1157.get(0);
        mod_1158.put(0, t);
    endrule
    rule rule_1514;
        ChannelMessage t;
        t <- mod_1153.get(3);
        mod_1154.put(0, t);
    endrule
    rule rule_1515;
        ChannelMessage t;
        t <- mod_1187.get(0);
        mod_1154.put(1, t);
    endrule
    rule rule_1516;
        ChannelMessage t;
        t <- mod_1172.get(0);
        mod_1160.put(1, t);
    endrule
    rule rule_1517;
        ChannelMessage t;
        t <- mod_1179.get(0);
        mod_1178.put(0, t);
    endrule
    rule rule_1518;
        ChannelMessage t;
        t <- mod_1183.get(0);
        mod_1182.put(1, t);
    endrule
    rule rule_1519;
        ChannelMessage t;
        t <- mod_1152.get(1);
        mod_1153.put(0, t);
    endrule
    rule rule_1520;
        ChannelMessage t;
        t <- mod_1154.get(0);
        mod_1187.put(0, t);
    endrule
    rule rule_1521;
        ChannelMessage t;
        t <- mod_1160.get(1);
        mod_1161.put(0, t);
    endrule
    rule rule_1522;
        ChannelMessage t;
        t <- mod_1171.get(0);
        mod_1170.put(0, t);
    endrule
    rule rule_1523;
        ChannelMessage t;
        t <- mod_1185.get(0);
        mod_1184.put(0, t);
    endrule
    rule rule_1524;
        ChannelMessage t;
        t <- mod_1178.get(0);
        mod_1176.put(0, t);
    endrule
    rule rule_1525;
        ChannelMessage t;
        t <- mod_1164.get(1);
        mod_1165.put(1, t);
    endrule
    rule rule_1526;
        ChannelMessage t;
        t <- mod_1151.get(0);
        mod_1152.put(0, t);
    endrule
    rule rule_1527;
        ChannelMessage t;
        t <- mod_1161.get(0);
        mod_1162.put(0, t);
    endrule
    rule rule_1528;
        ChannelMessage t;
        t <- mod_1174.get(0);
        mod_1173.put(0, t);
    endrule
    rule rule_1529;
        ChannelMessage t;
        t <- mod_1173.get(0);
        mod_1159.put(1, t);
    endrule
    rule rule_1530;
        ChannelMessage t;
        t <- mod_1175.get(0);
        mod_1174.put(0, t);
    endrule
    rule rule_1531;
        ChannelMessage t;
        t <- mod_1184.get(0);
        mod_1182.put(0, t);
    endrule
    rule rule_1532;
        ChannelMessage t;
        t <- mod_1154.get(1);
        mod_1155.put(0, t);
    endrule
    rule rule_1533;
        ChannelMessage t;
        t <- mod_1155.get(0);
        mod_1180.put(0, t);
    endrule
    rule rule_1534;
        ChannelMessage t;
        t <- mod_1168.get(1);
        mod_1161.put(1, t);
    endrule
    rule rule_1535;
        ChannelMessage t;
        t <- mod_1182.get(1);
        mod_1157.put(1, t);
    endrule
    rule rule_1536;
        ChannelMessage t;
        t <- mod_1188.get(1);
        mod_1152.put(1, t);
    endrule
    rule rule_1537;
        ChannelMessage t;
        t <- mod_1163.get(1);
        mod_1164.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1149.put(0, t);
        end
        if (i == 1) begin
            mod_1165.put(0, t);
        end
        if (i == 2) begin
            mod_1171.put(0, t);
        end
        if (i == 3) begin
            mod_1179.put(0, t);
        end
        if (i == 4) begin
            mod_1185.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_1153.get(0);
        end
        if (i == 1) begin
            t <- mod_1153.get(1);
        end
        if (i == 3) begin
            t <- mod_1153.get(2);
        end
        if (i == 2) begin
            t <- mod_1165.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6063 (Operation_IFC);
    Operation_IFC mod_1190_inner <- mkReshape(2, 64);
    Operation_IFC mod_1190 <- mkDebugOperation(mod_1190_inner, "mod_1190");
    Operation_IFC mod_1191_inner <- mkFlatten(1);
    Operation_IFC mod_1191 <- mkDebugOperation(mod_1191_inner, "mod_1191");
    Operation_IFC mod_1192_inner <- mkFlatten(2);
    Operation_IFC mod_1192 <- mkDebugOperation(mod_1192_inner, "mod_1192");
    Operation_IFC mod_1193_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1193 <- mkDebugOperation(mod_1193_inner, "mod_1193");
    Broadcast_IFC#(4) mod_1194_inner <- mkBroadcast(4);
    Operation_IFC mod_1194 <- mkDebugOperation(mod_1194_inner.op, "mod_1194");
    PMU_IFC mod_1195_bufferize <- mkPMU(2);
    Operation_IFC mod_1195_inner = mod_1195_bufferize.operation;
    Operation_IFC mod_1195 <- mkDebugOperation(mod_1195_inner, "mod_1195");
    Broadcast_IFC#(2) mod_1196_inner <- mkBroadcast(2);
    Operation_IFC mod_1196 <- mkDebugOperation(mod_1196_inner.op, "mod_1196");
    PMU_IFC mod_1197_bufferize <- mkPMU(1);
    Operation_IFC mod_1197_inner = mod_1197_bufferize.operation;
    Operation_IFC mod_1197 <- mkDebugOperation(mod_1197_inner, "mod_1197");
    Operation_IFC mod_1198_inner <- mkBinaryMap(1127, matmul_t_tile);
    Operation_IFC mod_1198 <- mkDebugOperation(mod_1198_inner, "mod_1198");
    Operation_IFC mod_1199_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1199 <- mkDebugOperation(mod_1199_inner, "mod_1199");
    Operation_IFC mod_1200_inner <- mkBinaryMap(1895, mul_tile);
    Operation_IFC mod_1200 <- mkDebugOperation(mod_1200_inner, "mod_1200");
    PMU_IFC mod_1201_bufferize <- mkPMU(1);
    Operation_IFC mod_1201_inner = mod_1201_bufferize.operation;
    Operation_IFC mod_1201 <- mkDebugOperation(mod_1201_inner, "mod_1201");
    Operation_IFC mod_1202_inner <- mkBinaryMap(2505, matmul_t_tile);
    Operation_IFC mod_1202 <- mkDebugOperation(mod_1202_inner, "mod_1202");
    Operation_IFC mod_1203_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1203 <- mkDebugOperation(mod_1203_inner, "mod_1203");
    Operation_IFC mod_1204_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1204 <- mkDebugOperation(mod_1204_inner, "mod_1204");
    Operation_IFC mod_1205_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1205 <- mkDebugOperation(mod_1205_inner, "mod_1205");
    Operation_IFC mod_1206_inner <- mkBinaryMap(2794, mul_tile);
    Operation_IFC mod_1206 <- mkDebugOperation(mod_1206_inner, "mod_1206");
    PMU_IFC mod_1207_bufferize <- mkPMU(1);
    Operation_IFC mod_1207_inner = mod_1207_bufferize.operation;
    Operation_IFC mod_1207 <- mkDebugOperation(mod_1207_inner, "mod_1207");
    PMU_IFC mod_1208_bufferize <- mkPMU(2);
    Operation_IFC mod_1208_inner = mod_1208_bufferize.operation;
    Operation_IFC mod_1208 <- mkDebugOperation(mod_1208_inner, "mod_1208");
    PMU_IFC mod_1209_bufferize <- mkPMU(2);
    Operation_IFC mod_1209_inner = mod_1209_bufferize.operation;
    Operation_IFC mod_1209 <- mkDebugOperation(mod_1209_inner, "mod_1209");
    Operation_IFC mod_1210_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1210 <- mkDebugOperation(mod_1210_inner, "mod_1210");
    Operation_IFC mod_1211_inner <- mkFlatten(1);
    Operation_IFC mod_1211 <- mkDebugOperation(mod_1211_inner, "mod_1211");
    Operation_IFC mod_1212_inner <- mkFlatten(0);
    Operation_IFC mod_1212 <- mkDebugOperation(mod_1212_inner, "mod_1212");
    Operation_IFC mod_1213_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1213 <- mkDebugOperation(mod_1213_inner, "mod_1213");
    Operation_IFC mod_1214_inner <- mkUnaryMap(1767, silu_tile);
    Operation_IFC mod_1214 <- mkDebugOperation(mod_1214_inner, "mod_1214");
    Operation_IFC mod_1215_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1215 <- mkDebugOperation(mod_1215_inner, "mod_1215");
    Operation_IFC mod_1216_inner <- mkBinaryMap(1639, matmul_t_tile);
    Operation_IFC mod_1216 <- mkDebugOperation(mod_1216_inner, "mod_1216");
    PMU_IFC mod_1217_bufferize <- mkPMU(2);
    Operation_IFC mod_1217_inner = mod_1217_bufferize.operation;
    Operation_IFC mod_1217 <- mkDebugOperation(mod_1217_inner, "mod_1217");
    Operation_IFC mod_1218_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1218 <- mkDebugOperation(mod_1218_inner, "mod_1218");
    Operation_IFC mod_1219_inner <- mkFlatten(1);
    Operation_IFC mod_1219 <- mkDebugOperation(mod_1219_inner, "mod_1219");
    Operation_IFC mod_1220_inner <- mkFlatten(0);
    Operation_IFC mod_1220 <- mkDebugOperation(mod_1220_inner, "mod_1220");
    PMU_IFC mod_1221_bufferize <- mkPMU(1);
    Operation_IFC mod_1221_inner = mod_1221_bufferize.operation;
    Operation_IFC mod_1221 <- mkDebugOperation(mod_1221_inner, "mod_1221");
    Operation_IFC mod_1222_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1222 <- mkDebugOperation(mod_1222_inner, "mod_1222");
    PMU_IFC mod_1223_bufferize <- mkPMU(2);
    Operation_IFC mod_1223_inner = mod_1223_bufferize.operation;
    Operation_IFC mod_1223 <- mkDebugOperation(mod_1223_inner, "mod_1223");
    Operation_IFC mod_1224_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1224 <- mkDebugOperation(mod_1224_inner, "mod_1224");
    Operation_IFC mod_1225_inner <- mkFlatten(1);
    Operation_IFC mod_1225 <- mkDebugOperation(mod_1225_inner, "mod_1225");
    Operation_IFC mod_1226_inner <- mkFlatten(0);
    Operation_IFC mod_1226 <- mkDebugOperation(mod_1226_inner, "mod_1226");
    Operation_IFC mod_1227_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1227 <- mkDebugOperation(mod_1227_inner, "mod_1227");
    Operation_IFC mod_1228_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1228 <- mkDebugOperation(mod_1228_inner, "mod_1228");
    PMU_IFC mod_1229_bufferize <- mkPMU(2);
    Operation_IFC mod_1229_inner = mod_1229_bufferize.operation;
    Operation_IFC mod_1229 <- mkDebugOperation(mod_1229_inner, "mod_1229");
    rule rule_1538;
        ChannelMessage t;
        t <- mod_1221.get(1);
        mod_1216.put(0, t);
    endrule
    rule rule_1539;
        ChannelMessage t;
        t <- mod_1225.get(0);
        mod_1223.put(0, t);
    endrule
    rule rule_1540;
        ChannelMessage t;
        t <- mod_1207.get(0);
        mod_1207.put(1, t);
    endrule
    rule rule_1541;
        ChannelMessage t;
        t <- mod_1227.get(0);
        mod_1197.put(1, t);
    endrule
    rule rule_1542;
        ChannelMessage t;
        t <- mod_1193.get(1);
        mod_1194.put(0, t);
    endrule
    rule rule_1543;
        ChannelMessage t;
        t <- mod_1222.get(0);
        mod_1221.put(1, t);
    endrule
    rule rule_1544;
        ChannelMessage t;
        t <- mod_1220.get(0);
        mod_1219.put(0, t);
    endrule
    rule rule_1545;
        ChannelMessage t;
        t <- mod_1221.get(0);
        mod_1222.put(0, t);
    endrule
    rule rule_1546;
        ChannelMessage t;
        t <- mod_1215.get(0);
        mod_1214.put(0, t);
    endrule
    rule rule_1547;
        ChannelMessage t;
        t <- mod_1195.get(1);
        mod_1196.put(0, t);
    endrule
    rule rule_1548;
        ChannelMessage t;
        t <- mod_1210.get(0);
        mod_1209.put(1, t);
    endrule
    rule rule_1549;
        ChannelMessage t;
        t <- mod_1205.get(1);
        mod_1206.put(1, t);
    endrule
    rule rule_1550;
        ChannelMessage t;
        t <- mod_1217.get(1);
        mod_1216.put(1, t);
    endrule
    rule rule_1551;
        ChannelMessage t;
        t <- mod_1213.get(0);
        mod_1201.put(1, t);
    endrule
    rule rule_1552;
        ChannelMessage t;
        t <- mod_1204.get(1);
        mod_1205.put(0, t);
    endrule
    rule rule_1553;
        ChannelMessage t;
        t <- mod_1228.get(0);
        mod_1195.put(1, t);
    endrule
    rule rule_1554;
        ChannelMessage t;
        t <- mod_1201.get(0);
        mod_1213.put(0, t);
    endrule
    rule rule_1555;
        ChannelMessage t;
        t <- mod_1209.get(1);
        mod_1202.put(1, t);
    endrule
    rule rule_1556;
        ChannelMessage t;
        t <- mod_1199.get(0);
        mod_1200.put(0, t);
    endrule
    rule rule_1557;
        ChannelMessage t;
        t <- mod_1219.get(0);
        mod_1217.put(0, t);
    endrule
    rule rule_1558;
        ChannelMessage t;
        t <- mod_1194.get(3);
        mod_1195.put(0, t);
    endrule
    rule rule_1559;
        ChannelMessage t;
        t <- mod_1201.get(1);
        mod_1202.put(0, t);
    endrule
    rule rule_1560;
        ChannelMessage t;
        t <- mod_1197.get(1);
        mod_1198.put(0, t);
    endrule
    rule rule_1561;
        ChannelMessage t;
        t <- mod_1209.get(0);
        mod_1210.put(0, t);
    endrule
    rule rule_1562;
        ChannelMessage t;
        t <- mod_1229.get(1);
        mod_1193.put(1, t);
    endrule
    rule rule_1563;
        ChannelMessage t;
        t <- mod_1202.get(0);
        mod_1203.put(0, t);
    endrule
    rule rule_1564;
        ChannelMessage t;
        t <- mod_1190.get(0);
        mod_1191.put(0, t);
    endrule
    rule rule_1565;
        ChannelMessage t;
        t <- mod_1226.get(0);
        mod_1225.put(0, t);
    endrule
    rule rule_1566;
        ChannelMessage t;
        t <- mod_1208.get(1);
        mod_1204.put(1, t);
    endrule
    rule rule_1567;
        ChannelMessage t;
        t <- mod_1192.get(0);
        mod_1193.put(0, t);
    endrule
    rule rule_1568;
        ChannelMessage t;
        t <- mod_1200.get(0);
        mod_1201.put(0, t);
    endrule
    rule rule_1569;
        ChannelMessage t;
        t <- mod_1211.get(0);
        mod_1209.put(0, t);
    endrule
    rule rule_1570;
        ChannelMessage t;
        t <- mod_1205.get(0);
        mod_1207.put(0, t);
    endrule
    rule rule_1571;
        ChannelMessage t;
        t <- mod_1197.get(0);
        mod_1227.put(0, t);
    endrule
    rule rule_1572;
        ChannelMessage t;
        t <- mod_1203.get(0);
        mod_1204.put(0, t);
    endrule
    rule rule_1573;
        ChannelMessage t;
        t <- mod_1212.get(0);
        mod_1211.put(0, t);
    endrule
    rule rule_1574;
        ChannelMessage t;
        t <- mod_1204.get(0);
        mod_1208.put(0, t);
    endrule
    rule rule_1575;
        ChannelMessage t;
        t <- mod_1216.get(0);
        mod_1215.put(0, t);
    endrule
    rule rule_1576;
        ChannelMessage t;
        t <- mod_1196.get(0);
        mod_1221.put(0, t);
    endrule
    rule rule_1577;
        ChannelMessage t;
        t <- mod_1229.get(0);
        mod_1229.put(1, t);
    endrule
    rule rule_1578;
        ChannelMessage t;
        t <- mod_1217.get(0);
        mod_1218.put(0, t);
    endrule
    rule rule_1579;
        ChannelMessage t;
        t <- mod_1223.get(1);
        mod_1198.put(1, t);
    endrule
    rule rule_1580;
        ChannelMessage t;
        t <- mod_1195.get(0);
        mod_1228.put(0, t);
    endrule
    rule rule_1581;
        ChannelMessage t;
        t <- mod_1198.get(0);
        mod_1199.put(0, t);
    endrule
    rule rule_1582;
        ChannelMessage t;
        t <- mod_1207.get(1);
        mod_1205.put(1, t);
    endrule
    rule rule_1583;
        ChannelMessage t;
        t <- mod_1218.get(0);
        mod_1217.put(1, t);
    endrule
    rule rule_1584;
        ChannelMessage t;
        t <- mod_1196.get(1);
        mod_1197.put(0, t);
    endrule
    rule rule_1585;
        ChannelMessage t;
        t <- mod_1193.get(0);
        mod_1229.put(0, t);
    endrule
    rule rule_1586;
        ChannelMessage t;
        t <- mod_1214.get(0);
        mod_1200.put(1, t);
    endrule
    rule rule_1587;
        ChannelMessage t;
        t <- mod_1224.get(0);
        mod_1223.put(1, t);
    endrule
    rule rule_1588;
        ChannelMessage t;
        t <- mod_1191.get(0);
        mod_1192.put(0, t);
    endrule
    rule rule_1589;
        ChannelMessage t;
        t <- mod_1208.get(0);
        mod_1208.put(1, t);
    endrule
    rule rule_1590;
        ChannelMessage t;
        t <- mod_1223.get(0);
        mod_1224.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1190.put(0, t);
        end
        if (i == 1) begin
            mod_1206.put(0, t);
        end
        if (i == 2) begin
            mod_1212.put(0, t);
        end
        if (i == 3) begin
            mod_1220.put(0, t);
        end
        if (i == 4) begin
            mod_1226.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_1194.get(0);
        end
        if (i == 0) begin
            t <- mod_1194.get(1);
        end
        if (i == 2) begin
            t <- mod_1194.get(2);
        end
        if (i == 3) begin
            t <- mod_1206.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6064 (Operation_IFC);
    Operation_IFC mod_1231_inner <- mkReshape(2, 64);
    Operation_IFC mod_1231 <- mkDebugOperation(mod_1231_inner, "mod_1231");
    Operation_IFC mod_1232_inner <- mkFlatten(1);
    Operation_IFC mod_1232 <- mkDebugOperation(mod_1232_inner, "mod_1232");
    Operation_IFC mod_1233_inner <- mkFlatten(2);
    Operation_IFC mod_1233 <- mkDebugOperation(mod_1233_inner, "mod_1233");
    Operation_IFC mod_1234_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1234 <- mkDebugOperation(mod_1234_inner, "mod_1234");
    Broadcast_IFC#(4) mod_1235_inner <- mkBroadcast(4);
    Operation_IFC mod_1235 <- mkDebugOperation(mod_1235_inner.op, "mod_1235");
    PMU_IFC mod_1236_bufferize <- mkPMU(2);
    Operation_IFC mod_1236_inner = mod_1236_bufferize.operation;
    Operation_IFC mod_1236 <- mkDebugOperation(mod_1236_inner, "mod_1236");
    Broadcast_IFC#(2) mod_1237_inner <- mkBroadcast(2);
    Operation_IFC mod_1237 <- mkDebugOperation(mod_1237_inner.op, "mod_1237");
    PMU_IFC mod_1238_bufferize <- mkPMU(1);
    Operation_IFC mod_1238_inner = mod_1238_bufferize.operation;
    Operation_IFC mod_1238 <- mkDebugOperation(mod_1238_inner, "mod_1238");
    Operation_IFC mod_1239_inner <- mkBinaryMap(1126, matmul_t_tile);
    Operation_IFC mod_1239 <- mkDebugOperation(mod_1239_inner, "mod_1239");
    Operation_IFC mod_1240_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1240 <- mkDebugOperation(mod_1240_inner, "mod_1240");
    Operation_IFC mod_1241_inner <- mkBinaryMap(1894, mul_tile);
    Operation_IFC mod_1241 <- mkDebugOperation(mod_1241_inner, "mod_1241");
    PMU_IFC mod_1242_bufferize <- mkPMU(1);
    Operation_IFC mod_1242_inner = mod_1242_bufferize.operation;
    Operation_IFC mod_1242 <- mkDebugOperation(mod_1242_inner, "mod_1242");
    Operation_IFC mod_1243_inner <- mkBinaryMap(2503, matmul_t_tile);
    Operation_IFC mod_1243 <- mkDebugOperation(mod_1243_inner, "mod_1243");
    Operation_IFC mod_1244_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1244 <- mkDebugOperation(mod_1244_inner, "mod_1244");
    Operation_IFC mod_1245_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1245 <- mkDebugOperation(mod_1245_inner, "mod_1245");
    Operation_IFC mod_1246_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1246 <- mkDebugOperation(mod_1246_inner, "mod_1246");
    Operation_IFC mod_1247_inner <- mkBinaryMap(2793, mul_tile);
    Operation_IFC mod_1247 <- mkDebugOperation(mod_1247_inner, "mod_1247");
    PMU_IFC mod_1248_bufferize <- mkPMU(1);
    Operation_IFC mod_1248_inner = mod_1248_bufferize.operation;
    Operation_IFC mod_1248 <- mkDebugOperation(mod_1248_inner, "mod_1248");
    PMU_IFC mod_1249_bufferize <- mkPMU(2);
    Operation_IFC mod_1249_inner = mod_1249_bufferize.operation;
    Operation_IFC mod_1249 <- mkDebugOperation(mod_1249_inner, "mod_1249");
    PMU_IFC mod_1250_bufferize <- mkPMU(2);
    Operation_IFC mod_1250_inner = mod_1250_bufferize.operation;
    Operation_IFC mod_1250 <- mkDebugOperation(mod_1250_inner, "mod_1250");
    Operation_IFC mod_1251_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1251 <- mkDebugOperation(mod_1251_inner, "mod_1251");
    Operation_IFC mod_1252_inner <- mkFlatten(1);
    Operation_IFC mod_1252 <- mkDebugOperation(mod_1252_inner, "mod_1252");
    Operation_IFC mod_1253_inner <- mkFlatten(0);
    Operation_IFC mod_1253 <- mkDebugOperation(mod_1253_inner, "mod_1253");
    Operation_IFC mod_1254_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1254 <- mkDebugOperation(mod_1254_inner, "mod_1254");
    Operation_IFC mod_1255_inner <- mkUnaryMap(1766, silu_tile);
    Operation_IFC mod_1255 <- mkDebugOperation(mod_1255_inner, "mod_1255");
    Operation_IFC mod_1256_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1256 <- mkDebugOperation(mod_1256_inner, "mod_1256");
    Operation_IFC mod_1257_inner <- mkBinaryMap(1638, matmul_t_tile);
    Operation_IFC mod_1257 <- mkDebugOperation(mod_1257_inner, "mod_1257");
    PMU_IFC mod_1258_bufferize <- mkPMU(2);
    Operation_IFC mod_1258_inner = mod_1258_bufferize.operation;
    Operation_IFC mod_1258 <- mkDebugOperation(mod_1258_inner, "mod_1258");
    Operation_IFC mod_1259_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1259 <- mkDebugOperation(mod_1259_inner, "mod_1259");
    Operation_IFC mod_1260_inner <- mkFlatten(1);
    Operation_IFC mod_1260 <- mkDebugOperation(mod_1260_inner, "mod_1260");
    Operation_IFC mod_1261_inner <- mkFlatten(0);
    Operation_IFC mod_1261 <- mkDebugOperation(mod_1261_inner, "mod_1261");
    PMU_IFC mod_1262_bufferize <- mkPMU(1);
    Operation_IFC mod_1262_inner = mod_1262_bufferize.operation;
    Operation_IFC mod_1262 <- mkDebugOperation(mod_1262_inner, "mod_1262");
    Operation_IFC mod_1263_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1263 <- mkDebugOperation(mod_1263_inner, "mod_1263");
    PMU_IFC mod_1264_bufferize <- mkPMU(2);
    Operation_IFC mod_1264_inner = mod_1264_bufferize.operation;
    Operation_IFC mod_1264 <- mkDebugOperation(mod_1264_inner, "mod_1264");
    Operation_IFC mod_1265_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1265 <- mkDebugOperation(mod_1265_inner, "mod_1265");
    Operation_IFC mod_1266_inner <- mkFlatten(1);
    Operation_IFC mod_1266 <- mkDebugOperation(mod_1266_inner, "mod_1266");
    Operation_IFC mod_1267_inner <- mkFlatten(0);
    Operation_IFC mod_1267 <- mkDebugOperation(mod_1267_inner, "mod_1267");
    Operation_IFC mod_1268_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1268 <- mkDebugOperation(mod_1268_inner, "mod_1268");
    Operation_IFC mod_1269_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1269 <- mkDebugOperation(mod_1269_inner, "mod_1269");
    PMU_IFC mod_1270_bufferize <- mkPMU(2);
    Operation_IFC mod_1270_inner = mod_1270_bufferize.operation;
    Operation_IFC mod_1270 <- mkDebugOperation(mod_1270_inner, "mod_1270");
    rule rule_1591;
        ChannelMessage t;
        t <- mod_1252.get(0);
        mod_1250.put(0, t);
    endrule
    rule rule_1592;
        ChannelMessage t;
        t <- mod_1231.get(0);
        mod_1232.put(0, t);
    endrule
    rule rule_1593;
        ChannelMessage t;
        t <- mod_1237.get(0);
        mod_1262.put(0, t);
    endrule
    rule rule_1594;
        ChannelMessage t;
        t <- mod_1246.get(0);
        mod_1248.put(0, t);
    endrule
    rule rule_1595;
        ChannelMessage t;
        t <- mod_1256.get(0);
        mod_1255.put(0, t);
    endrule
    rule rule_1596;
        ChannelMessage t;
        t <- mod_1234.get(0);
        mod_1270.put(0, t);
    endrule
    rule rule_1597;
        ChannelMessage t;
        t <- mod_1246.get(1);
        mod_1247.put(1, t);
    endrule
    rule rule_1598;
        ChannelMessage t;
        t <- mod_1250.get(1);
        mod_1243.put(1, t);
    endrule
    rule rule_1599;
        ChannelMessage t;
        t <- mod_1242.get(1);
        mod_1243.put(0, t);
    endrule
    rule rule_1600;
        ChannelMessage t;
        t <- mod_1258.get(0);
        mod_1259.put(0, t);
    endrule
    rule rule_1601;
        ChannelMessage t;
        t <- mod_1265.get(0);
        mod_1264.put(1, t);
    endrule
    rule rule_1602;
        ChannelMessage t;
        t <- mod_1245.get(1);
        mod_1246.put(0, t);
    endrule
    rule rule_1603;
        ChannelMessage t;
        t <- mod_1248.get(1);
        mod_1246.put(1, t);
    endrule
    rule rule_1604;
        ChannelMessage t;
        t <- mod_1245.get(0);
        mod_1249.put(0, t);
    endrule
    rule rule_1605;
        ChannelMessage t;
        t <- mod_1249.get(1);
        mod_1245.put(1, t);
    endrule
    rule rule_1606;
        ChannelMessage t;
        t <- mod_1236.get(0);
        mod_1269.put(0, t);
    endrule
    rule rule_1607;
        ChannelMessage t;
        t <- mod_1264.get(0);
        mod_1265.put(0, t);
    endrule
    rule rule_1608;
        ChannelMessage t;
        t <- mod_1270.get(1);
        mod_1234.put(1, t);
    endrule
    rule rule_1609;
        ChannelMessage t;
        t <- mod_1262.get(0);
        mod_1263.put(0, t);
    endrule
    rule rule_1610;
        ChannelMessage t;
        t <- mod_1238.get(0);
        mod_1268.put(0, t);
    endrule
    rule rule_1611;
        ChannelMessage t;
        t <- mod_1250.get(0);
        mod_1251.put(0, t);
    endrule
    rule rule_1612;
        ChannelMessage t;
        t <- mod_1253.get(0);
        mod_1252.put(0, t);
    endrule
    rule rule_1613;
        ChannelMessage t;
        t <- mod_1263.get(0);
        mod_1262.put(1, t);
    endrule
    rule rule_1614;
        ChannelMessage t;
        t <- mod_1268.get(0);
        mod_1238.put(1, t);
    endrule
    rule rule_1615;
        ChannelMessage t;
        t <- mod_1269.get(0);
        mod_1236.put(1, t);
    endrule
    rule rule_1616;
        ChannelMessage t;
        t <- mod_1258.get(1);
        mod_1257.put(1, t);
    endrule
    rule rule_1617;
        ChannelMessage t;
        t <- mod_1242.get(0);
        mod_1254.put(0, t);
    endrule
    rule rule_1618;
        ChannelMessage t;
        t <- mod_1254.get(0);
        mod_1242.put(1, t);
    endrule
    rule rule_1619;
        ChannelMessage t;
        t <- mod_1233.get(0);
        mod_1234.put(0, t);
    endrule
    rule rule_1620;
        ChannelMessage t;
        t <- mod_1236.get(1);
        mod_1237.put(0, t);
    endrule
    rule rule_1621;
        ChannelMessage t;
        t <- mod_1255.get(0);
        mod_1241.put(1, t);
    endrule
    rule rule_1622;
        ChannelMessage t;
        t <- mod_1248.get(0);
        mod_1248.put(1, t);
    endrule
    rule rule_1623;
        ChannelMessage t;
        t <- mod_1259.get(0);
        mod_1258.put(1, t);
    endrule
    rule rule_1624;
        ChannelMessage t;
        t <- mod_1270.get(0);
        mod_1270.put(1, t);
    endrule
    rule rule_1625;
        ChannelMessage t;
        t <- mod_1239.get(0);
        mod_1240.put(0, t);
    endrule
    rule rule_1626;
        ChannelMessage t;
        t <- mod_1232.get(0);
        mod_1233.put(0, t);
    endrule
    rule rule_1627;
        ChannelMessage t;
        t <- mod_1267.get(0);
        mod_1266.put(0, t);
    endrule
    rule rule_1628;
        ChannelMessage t;
        t <- mod_1243.get(0);
        mod_1244.put(0, t);
    endrule
    rule rule_1629;
        ChannelMessage t;
        t <- mod_1235.get(3);
        mod_1236.put(0, t);
    endrule
    rule rule_1630;
        ChannelMessage t;
        t <- mod_1251.get(0);
        mod_1250.put(1, t);
    endrule
    rule rule_1631;
        ChannelMessage t;
        t <- mod_1260.get(0);
        mod_1258.put(0, t);
    endrule
    rule rule_1632;
        ChannelMessage t;
        t <- mod_1261.get(0);
        mod_1260.put(0, t);
    endrule
    rule rule_1633;
        ChannelMessage t;
        t <- mod_1234.get(1);
        mod_1235.put(0, t);
    endrule
    rule rule_1634;
        ChannelMessage t;
        t <- mod_1240.get(0);
        mod_1241.put(0, t);
    endrule
    rule rule_1635;
        ChannelMessage t;
        t <- mod_1241.get(0);
        mod_1242.put(0, t);
    endrule
    rule rule_1636;
        ChannelMessage t;
        t <- mod_1249.get(0);
        mod_1249.put(1, t);
    endrule
    rule rule_1637;
        ChannelMessage t;
        t <- mod_1262.get(1);
        mod_1257.put(0, t);
    endrule
    rule rule_1638;
        ChannelMessage t;
        t <- mod_1244.get(0);
        mod_1245.put(0, t);
    endrule
    rule rule_1639;
        ChannelMessage t;
        t <- mod_1238.get(1);
        mod_1239.put(0, t);
    endrule
    rule rule_1640;
        ChannelMessage t;
        t <- mod_1257.get(0);
        mod_1256.put(0, t);
    endrule
    rule rule_1641;
        ChannelMessage t;
        t <- mod_1266.get(0);
        mod_1264.put(0, t);
    endrule
    rule rule_1642;
        ChannelMessage t;
        t <- mod_1237.get(1);
        mod_1238.put(0, t);
    endrule
    rule rule_1643;
        ChannelMessage t;
        t <- mod_1264.get(1);
        mod_1239.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1231.put(0, t);
        end
        if (i == 1) begin
            mod_1247.put(0, t);
        end
        if (i == 2) begin
            mod_1253.put(0, t);
        end
        if (i == 3) begin
            mod_1261.put(0, t);
        end
        if (i == 4) begin
            mod_1267.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_1235.get(0);
        end
        if (i == 1) begin
            t <- mod_1235.get(1);
        end
        if (i == 0) begin
            t <- mod_1235.get(2);
        end
        if (i == 2) begin
            t <- mod_1247.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6065 (Operation_IFC);
    Operation_IFC mod_1272_inner <- mkReshape(2, 64);
    Operation_IFC mod_1272 <- mkDebugOperation(mod_1272_inner, "mod_1272");
    Operation_IFC mod_1273_inner <- mkFlatten(1);
    Operation_IFC mod_1273 <- mkDebugOperation(mod_1273_inner, "mod_1273");
    Operation_IFC mod_1274_inner <- mkFlatten(2);
    Operation_IFC mod_1274 <- mkDebugOperation(mod_1274_inner, "mod_1274");
    Operation_IFC mod_1275_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1275 <- mkDebugOperation(mod_1275_inner, "mod_1275");
    Broadcast_IFC#(4) mod_1276_inner <- mkBroadcast(4);
    Operation_IFC mod_1276 <- mkDebugOperation(mod_1276_inner.op, "mod_1276");
    PMU_IFC mod_1277_bufferize <- mkPMU(2);
    Operation_IFC mod_1277_inner = mod_1277_bufferize.operation;
    Operation_IFC mod_1277 <- mkDebugOperation(mod_1277_inner, "mod_1277");
    Broadcast_IFC#(2) mod_1278_inner <- mkBroadcast(2);
    Operation_IFC mod_1278 <- mkDebugOperation(mod_1278_inner.op, "mod_1278");
    PMU_IFC mod_1279_bufferize <- mkPMU(1);
    Operation_IFC mod_1279_inner = mod_1279_bufferize.operation;
    Operation_IFC mod_1279 <- mkDebugOperation(mod_1279_inner, "mod_1279");
    Operation_IFC mod_1280_inner <- mkBinaryMap(1125, matmul_t_tile);
    Operation_IFC mod_1280 <- mkDebugOperation(mod_1280_inner, "mod_1280");
    Operation_IFC mod_1281_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1281 <- mkDebugOperation(mod_1281_inner, "mod_1281");
    Operation_IFC mod_1282_inner <- mkBinaryMap(1893, mul_tile);
    Operation_IFC mod_1282 <- mkDebugOperation(mod_1282_inner, "mod_1282");
    PMU_IFC mod_1283_bufferize <- mkPMU(1);
    Operation_IFC mod_1283_inner = mod_1283_bufferize.operation;
    Operation_IFC mod_1283 <- mkDebugOperation(mod_1283_inner, "mod_1283");
    Operation_IFC mod_1284_inner <- mkBinaryMap(2501, matmul_t_tile);
    Operation_IFC mod_1284 <- mkDebugOperation(mod_1284_inner, "mod_1284");
    Operation_IFC mod_1285_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1285 <- mkDebugOperation(mod_1285_inner, "mod_1285");
    Operation_IFC mod_1286_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1286 <- mkDebugOperation(mod_1286_inner, "mod_1286");
    Operation_IFC mod_1287_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1287 <- mkDebugOperation(mod_1287_inner, "mod_1287");
    Operation_IFC mod_1288_inner <- mkBinaryMap(2792, mul_tile);
    Operation_IFC mod_1288 <- mkDebugOperation(mod_1288_inner, "mod_1288");
    PMU_IFC mod_1289_bufferize <- mkPMU(1);
    Operation_IFC mod_1289_inner = mod_1289_bufferize.operation;
    Operation_IFC mod_1289 <- mkDebugOperation(mod_1289_inner, "mod_1289");
    PMU_IFC mod_1290_bufferize <- mkPMU(2);
    Operation_IFC mod_1290_inner = mod_1290_bufferize.operation;
    Operation_IFC mod_1290 <- mkDebugOperation(mod_1290_inner, "mod_1290");
    PMU_IFC mod_1291_bufferize <- mkPMU(2);
    Operation_IFC mod_1291_inner = mod_1291_bufferize.operation;
    Operation_IFC mod_1291 <- mkDebugOperation(mod_1291_inner, "mod_1291");
    Operation_IFC mod_1292_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1292 <- mkDebugOperation(mod_1292_inner, "mod_1292");
    Operation_IFC mod_1293_inner <- mkFlatten(1);
    Operation_IFC mod_1293 <- mkDebugOperation(mod_1293_inner, "mod_1293");
    Operation_IFC mod_1294_inner <- mkFlatten(0);
    Operation_IFC mod_1294 <- mkDebugOperation(mod_1294_inner, "mod_1294");
    Operation_IFC mod_1295_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1295 <- mkDebugOperation(mod_1295_inner, "mod_1295");
    Operation_IFC mod_1296_inner <- mkUnaryMap(1765, silu_tile);
    Operation_IFC mod_1296 <- mkDebugOperation(mod_1296_inner, "mod_1296");
    Operation_IFC mod_1297_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1297 <- mkDebugOperation(mod_1297_inner, "mod_1297");
    Operation_IFC mod_1298_inner <- mkBinaryMap(1637, matmul_t_tile);
    Operation_IFC mod_1298 <- mkDebugOperation(mod_1298_inner, "mod_1298");
    PMU_IFC mod_1299_bufferize <- mkPMU(2);
    Operation_IFC mod_1299_inner = mod_1299_bufferize.operation;
    Operation_IFC mod_1299 <- mkDebugOperation(mod_1299_inner, "mod_1299");
    Operation_IFC mod_1300_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1300 <- mkDebugOperation(mod_1300_inner, "mod_1300");
    Operation_IFC mod_1301_inner <- mkFlatten(1);
    Operation_IFC mod_1301 <- mkDebugOperation(mod_1301_inner, "mod_1301");
    Operation_IFC mod_1302_inner <- mkFlatten(0);
    Operation_IFC mod_1302 <- mkDebugOperation(mod_1302_inner, "mod_1302");
    PMU_IFC mod_1303_bufferize <- mkPMU(1);
    Operation_IFC mod_1303_inner = mod_1303_bufferize.operation;
    Operation_IFC mod_1303 <- mkDebugOperation(mod_1303_inner, "mod_1303");
    Operation_IFC mod_1304_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1304 <- mkDebugOperation(mod_1304_inner, "mod_1304");
    PMU_IFC mod_1305_bufferize <- mkPMU(2);
    Operation_IFC mod_1305_inner = mod_1305_bufferize.operation;
    Operation_IFC mod_1305 <- mkDebugOperation(mod_1305_inner, "mod_1305");
    Operation_IFC mod_1306_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1306 <- mkDebugOperation(mod_1306_inner, "mod_1306");
    Operation_IFC mod_1307_inner <- mkFlatten(1);
    Operation_IFC mod_1307 <- mkDebugOperation(mod_1307_inner, "mod_1307");
    Operation_IFC mod_1308_inner <- mkFlatten(0);
    Operation_IFC mod_1308 <- mkDebugOperation(mod_1308_inner, "mod_1308");
    Operation_IFC mod_1309_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1309 <- mkDebugOperation(mod_1309_inner, "mod_1309");
    Operation_IFC mod_1310_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1310 <- mkDebugOperation(mod_1310_inner, "mod_1310");
    PMU_IFC mod_1311_bufferize <- mkPMU(2);
    Operation_IFC mod_1311_inner = mod_1311_bufferize.operation;
    Operation_IFC mod_1311 <- mkDebugOperation(mod_1311_inner, "mod_1311");
    rule rule_1644;
        ChannelMessage t;
        t <- mod_1273.get(0);
        mod_1274.put(0, t);
    endrule
    rule rule_1645;
        ChannelMessage t;
        t <- mod_1293.get(0);
        mod_1291.put(0, t);
    endrule
    rule rule_1646;
        ChannelMessage t;
        t <- mod_1300.get(0);
        mod_1299.put(1, t);
    endrule
    rule rule_1647;
        ChannelMessage t;
        t <- mod_1303.get(1);
        mod_1298.put(0, t);
    endrule
    rule rule_1648;
        ChannelMessage t;
        t <- mod_1281.get(0);
        mod_1282.put(0, t);
    endrule
    rule rule_1649;
        ChannelMessage t;
        t <- mod_1290.get(0);
        mod_1290.put(1, t);
    endrule
    rule rule_1650;
        ChannelMessage t;
        t <- mod_1292.get(0);
        mod_1291.put(1, t);
    endrule
    rule rule_1651;
        ChannelMessage t;
        t <- mod_1278.get(0);
        mod_1303.put(0, t);
    endrule
    rule rule_1652;
        ChannelMessage t;
        t <- mod_1303.get(0);
        mod_1304.put(0, t);
    endrule
    rule rule_1653;
        ChannelMessage t;
        t <- mod_1297.get(0);
        mod_1296.put(0, t);
    endrule
    rule rule_1654;
        ChannelMessage t;
        t <- mod_1280.get(0);
        mod_1281.put(0, t);
    endrule
    rule rule_1655;
        ChannelMessage t;
        t <- mod_1310.get(0);
        mod_1277.put(1, t);
    endrule
    rule rule_1656;
        ChannelMessage t;
        t <- mod_1277.get(0);
        mod_1310.put(0, t);
    endrule
    rule rule_1657;
        ChannelMessage t;
        t <- mod_1276.get(3);
        mod_1277.put(0, t);
    endrule
    rule rule_1658;
        ChannelMessage t;
        t <- mod_1279.get(1);
        mod_1280.put(0, t);
    endrule
    rule rule_1659;
        ChannelMessage t;
        t <- mod_1275.get(1);
        mod_1276.put(0, t);
    endrule
    rule rule_1660;
        ChannelMessage t;
        t <- mod_1289.get(1);
        mod_1287.put(1, t);
    endrule
    rule rule_1661;
        ChannelMessage t;
        t <- mod_1286.get(0);
        mod_1290.put(0, t);
    endrule
    rule rule_1662;
        ChannelMessage t;
        t <- mod_1274.get(0);
        mod_1275.put(0, t);
    endrule
    rule rule_1663;
        ChannelMessage t;
        t <- mod_1286.get(1);
        mod_1287.put(0, t);
    endrule
    rule rule_1664;
        ChannelMessage t;
        t <- mod_1272.get(0);
        mod_1273.put(0, t);
    endrule
    rule rule_1665;
        ChannelMessage t;
        t <- mod_1284.get(0);
        mod_1285.put(0, t);
    endrule
    rule rule_1666;
        ChannelMessage t;
        t <- mod_1307.get(0);
        mod_1305.put(0, t);
    endrule
    rule rule_1667;
        ChannelMessage t;
        t <- mod_1295.get(0);
        mod_1283.put(1, t);
    endrule
    rule rule_1668;
        ChannelMessage t;
        t <- mod_1287.get(0);
        mod_1289.put(0, t);
    endrule
    rule rule_1669;
        ChannelMessage t;
        t <- mod_1283.get(1);
        mod_1284.put(0, t);
    endrule
    rule rule_1670;
        ChannelMessage t;
        t <- mod_1304.get(0);
        mod_1303.put(1, t);
    endrule
    rule rule_1671;
        ChannelMessage t;
        t <- mod_1296.get(0);
        mod_1282.put(1, t);
    endrule
    rule rule_1672;
        ChannelMessage t;
        t <- mod_1301.get(0);
        mod_1299.put(0, t);
    endrule
    rule rule_1673;
        ChannelMessage t;
        t <- mod_1277.get(1);
        mod_1278.put(0, t);
    endrule
    rule rule_1674;
        ChannelMessage t;
        t <- mod_1299.get(1);
        mod_1298.put(1, t);
    endrule
    rule rule_1675;
        ChannelMessage t;
        t <- mod_1291.get(0);
        mod_1292.put(0, t);
    endrule
    rule rule_1676;
        ChannelMessage t;
        t <- mod_1287.get(1);
        mod_1288.put(1, t);
    endrule
    rule rule_1677;
        ChannelMessage t;
        t <- mod_1278.get(1);
        mod_1279.put(0, t);
    endrule
    rule rule_1678;
        ChannelMessage t;
        t <- mod_1302.get(0);
        mod_1301.put(0, t);
    endrule
    rule rule_1679;
        ChannelMessage t;
        t <- mod_1311.get(1);
        mod_1275.put(1, t);
    endrule
    rule rule_1680;
        ChannelMessage t;
        t <- mod_1309.get(0);
        mod_1279.put(1, t);
    endrule
    rule rule_1681;
        ChannelMessage t;
        t <- mod_1289.get(0);
        mod_1289.put(1, t);
    endrule
    rule rule_1682;
        ChannelMessage t;
        t <- mod_1279.get(0);
        mod_1309.put(0, t);
    endrule
    rule rule_1683;
        ChannelMessage t;
        t <- mod_1306.get(0);
        mod_1305.put(1, t);
    endrule
    rule rule_1684;
        ChannelMessage t;
        t <- mod_1305.get(0);
        mod_1306.put(0, t);
    endrule
    rule rule_1685;
        ChannelMessage t;
        t <- mod_1299.get(0);
        mod_1300.put(0, t);
    endrule
    rule rule_1686;
        ChannelMessage t;
        t <- mod_1275.get(0);
        mod_1311.put(0, t);
    endrule
    rule rule_1687;
        ChannelMessage t;
        t <- mod_1283.get(0);
        mod_1295.put(0, t);
    endrule
    rule rule_1688;
        ChannelMessage t;
        t <- mod_1305.get(1);
        mod_1280.put(1, t);
    endrule
    rule rule_1689;
        ChannelMessage t;
        t <- mod_1308.get(0);
        mod_1307.put(0, t);
    endrule
    rule rule_1690;
        ChannelMessage t;
        t <- mod_1298.get(0);
        mod_1297.put(0, t);
    endrule
    rule rule_1691;
        ChannelMessage t;
        t <- mod_1291.get(1);
        mod_1284.put(1, t);
    endrule
    rule rule_1692;
        ChannelMessage t;
        t <- mod_1282.get(0);
        mod_1283.put(0, t);
    endrule
    rule rule_1693;
        ChannelMessage t;
        t <- mod_1294.get(0);
        mod_1293.put(0, t);
    endrule
    rule rule_1694;
        ChannelMessage t;
        t <- mod_1290.get(1);
        mod_1286.put(1, t);
    endrule
    rule rule_1695;
        ChannelMessage t;
        t <- mod_1285.get(0);
        mod_1286.put(0, t);
    endrule
    rule rule_1696;
        ChannelMessage t;
        t <- mod_1311.get(0);
        mod_1311.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1272.put(0, t);
        end
        if (i == 1) begin
            mod_1288.put(0, t);
        end
        if (i == 2) begin
            mod_1294.put(0, t);
        end
        if (i == 3) begin
            mod_1302.put(0, t);
        end
        if (i == 4) begin
            mod_1308.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_1276.get(0);
        end
        if (i == 3) begin
            t <- mod_1276.get(1);
        end
        if (i == 1) begin
            t <- mod_1276.get(2);
        end
        if (i == 2) begin
            t <- mod_1288.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6066 (Operation_IFC);
    Operation_IFC mod_1313_inner <- mkReshape(2, 64);
    Operation_IFC mod_1313 <- mkDebugOperation(mod_1313_inner, "mod_1313");
    Operation_IFC mod_1314_inner <- mkFlatten(1);
    Operation_IFC mod_1314 <- mkDebugOperation(mod_1314_inner, "mod_1314");
    Operation_IFC mod_1315_inner <- mkFlatten(2);
    Operation_IFC mod_1315 <- mkDebugOperation(mod_1315_inner, "mod_1315");
    Operation_IFC mod_1316_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1316 <- mkDebugOperation(mod_1316_inner, "mod_1316");
    Broadcast_IFC#(4) mod_1317_inner <- mkBroadcast(4);
    Operation_IFC mod_1317 <- mkDebugOperation(mod_1317_inner.op, "mod_1317");
    PMU_IFC mod_1318_bufferize <- mkPMU(2);
    Operation_IFC mod_1318_inner = mod_1318_bufferize.operation;
    Operation_IFC mod_1318 <- mkDebugOperation(mod_1318_inner, "mod_1318");
    Broadcast_IFC#(2) mod_1319_inner <- mkBroadcast(2);
    Operation_IFC mod_1319 <- mkDebugOperation(mod_1319_inner.op, "mod_1319");
    PMU_IFC mod_1320_bufferize <- mkPMU(1);
    Operation_IFC mod_1320_inner = mod_1320_bufferize.operation;
    Operation_IFC mod_1320 <- mkDebugOperation(mod_1320_inner, "mod_1320");
    Operation_IFC mod_1321_inner <- mkBinaryMap(1124, matmul_t_tile);
    Operation_IFC mod_1321 <- mkDebugOperation(mod_1321_inner, "mod_1321");
    Operation_IFC mod_1322_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1322 <- mkDebugOperation(mod_1322_inner, "mod_1322");
    Operation_IFC mod_1323_inner <- mkBinaryMap(1892, mul_tile);
    Operation_IFC mod_1323 <- mkDebugOperation(mod_1323_inner, "mod_1323");
    PMU_IFC mod_1324_bufferize <- mkPMU(1);
    Operation_IFC mod_1324_inner = mod_1324_bufferize.operation;
    Operation_IFC mod_1324 <- mkDebugOperation(mod_1324_inner, "mod_1324");
    Operation_IFC mod_1325_inner <- mkBinaryMap(2499, matmul_t_tile);
    Operation_IFC mod_1325 <- mkDebugOperation(mod_1325_inner, "mod_1325");
    Operation_IFC mod_1326_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1326 <- mkDebugOperation(mod_1326_inner, "mod_1326");
    Operation_IFC mod_1327_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1327 <- mkDebugOperation(mod_1327_inner, "mod_1327");
    Operation_IFC mod_1328_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1328 <- mkDebugOperation(mod_1328_inner, "mod_1328");
    Operation_IFC mod_1329_inner <- mkBinaryMap(2791, mul_tile);
    Operation_IFC mod_1329 <- mkDebugOperation(mod_1329_inner, "mod_1329");
    PMU_IFC mod_1330_bufferize <- mkPMU(1);
    Operation_IFC mod_1330_inner = mod_1330_bufferize.operation;
    Operation_IFC mod_1330 <- mkDebugOperation(mod_1330_inner, "mod_1330");
    PMU_IFC mod_1331_bufferize <- mkPMU(2);
    Operation_IFC mod_1331_inner = mod_1331_bufferize.operation;
    Operation_IFC mod_1331 <- mkDebugOperation(mod_1331_inner, "mod_1331");
    PMU_IFC mod_1332_bufferize <- mkPMU(2);
    Operation_IFC mod_1332_inner = mod_1332_bufferize.operation;
    Operation_IFC mod_1332 <- mkDebugOperation(mod_1332_inner, "mod_1332");
    Operation_IFC mod_1333_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1333 <- mkDebugOperation(mod_1333_inner, "mod_1333");
    Operation_IFC mod_1334_inner <- mkFlatten(1);
    Operation_IFC mod_1334 <- mkDebugOperation(mod_1334_inner, "mod_1334");
    Operation_IFC mod_1335_inner <- mkFlatten(0);
    Operation_IFC mod_1335 <- mkDebugOperation(mod_1335_inner, "mod_1335");
    Operation_IFC mod_1336_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1336 <- mkDebugOperation(mod_1336_inner, "mod_1336");
    Operation_IFC mod_1337_inner <- mkUnaryMap(1764, silu_tile);
    Operation_IFC mod_1337 <- mkDebugOperation(mod_1337_inner, "mod_1337");
    Operation_IFC mod_1338_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1338 <- mkDebugOperation(mod_1338_inner, "mod_1338");
    Operation_IFC mod_1339_inner <- mkBinaryMap(1636, matmul_t_tile);
    Operation_IFC mod_1339 <- mkDebugOperation(mod_1339_inner, "mod_1339");
    PMU_IFC mod_1340_bufferize <- mkPMU(2);
    Operation_IFC mod_1340_inner = mod_1340_bufferize.operation;
    Operation_IFC mod_1340 <- mkDebugOperation(mod_1340_inner, "mod_1340");
    Operation_IFC mod_1341_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1341 <- mkDebugOperation(mod_1341_inner, "mod_1341");
    Operation_IFC mod_1342_inner <- mkFlatten(1);
    Operation_IFC mod_1342 <- mkDebugOperation(mod_1342_inner, "mod_1342");
    Operation_IFC mod_1343_inner <- mkFlatten(0);
    Operation_IFC mod_1343 <- mkDebugOperation(mod_1343_inner, "mod_1343");
    PMU_IFC mod_1344_bufferize <- mkPMU(1);
    Operation_IFC mod_1344_inner = mod_1344_bufferize.operation;
    Operation_IFC mod_1344 <- mkDebugOperation(mod_1344_inner, "mod_1344");
    Operation_IFC mod_1345_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1345 <- mkDebugOperation(mod_1345_inner, "mod_1345");
    PMU_IFC mod_1346_bufferize <- mkPMU(2);
    Operation_IFC mod_1346_inner = mod_1346_bufferize.operation;
    Operation_IFC mod_1346 <- mkDebugOperation(mod_1346_inner, "mod_1346");
    Operation_IFC mod_1347_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1347 <- mkDebugOperation(mod_1347_inner, "mod_1347");
    Operation_IFC mod_1348_inner <- mkFlatten(1);
    Operation_IFC mod_1348 <- mkDebugOperation(mod_1348_inner, "mod_1348");
    Operation_IFC mod_1349_inner <- mkFlatten(0);
    Operation_IFC mod_1349 <- mkDebugOperation(mod_1349_inner, "mod_1349");
    Operation_IFC mod_1350_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1350 <- mkDebugOperation(mod_1350_inner, "mod_1350");
    Operation_IFC mod_1351_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1351 <- mkDebugOperation(mod_1351_inner, "mod_1351");
    PMU_IFC mod_1352_bufferize <- mkPMU(2);
    Operation_IFC mod_1352_inner = mod_1352_bufferize.operation;
    Operation_IFC mod_1352 <- mkDebugOperation(mod_1352_inner, "mod_1352");
    rule rule_1697;
        ChannelMessage t;
        t <- mod_1333.get(0);
        mod_1332.put(1, t);
    endrule
    rule rule_1698;
        ChannelMessage t;
        t <- mod_1331.get(1);
        mod_1327.put(1, t);
    endrule
    rule rule_1699;
        ChannelMessage t;
        t <- mod_1336.get(0);
        mod_1324.put(1, t);
    endrule
    rule rule_1700;
        ChannelMessage t;
        t <- mod_1347.get(0);
        mod_1346.put(1, t);
    endrule
    rule rule_1701;
        ChannelMessage t;
        t <- mod_1324.get(1);
        mod_1325.put(0, t);
    endrule
    rule rule_1702;
        ChannelMessage t;
        t <- mod_1340.get(0);
        mod_1341.put(0, t);
    endrule
    rule rule_1703;
        ChannelMessage t;
        t <- mod_1344.get(0);
        mod_1345.put(0, t);
    endrule
    rule rule_1704;
        ChannelMessage t;
        t <- mod_1328.get(1);
        mod_1329.put(1, t);
    endrule
    rule rule_1705;
        ChannelMessage t;
        t <- mod_1327.get(0);
        mod_1331.put(0, t);
    endrule
    rule rule_1706;
        ChannelMessage t;
        t <- mod_1330.get(0);
        mod_1330.put(1, t);
    endrule
    rule rule_1707;
        ChannelMessage t;
        t <- mod_1346.get(0);
        mod_1347.put(0, t);
    endrule
    rule rule_1708;
        ChannelMessage t;
        t <- mod_1320.get(0);
        mod_1350.put(0, t);
    endrule
    rule rule_1709;
        ChannelMessage t;
        t <- mod_1323.get(0);
        mod_1324.put(0, t);
    endrule
    rule rule_1710;
        ChannelMessage t;
        t <- mod_1338.get(0);
        mod_1337.put(0, t);
    endrule
    rule rule_1711;
        ChannelMessage t;
        t <- mod_1318.get(1);
        mod_1319.put(0, t);
    endrule
    rule rule_1712;
        ChannelMessage t;
        t <- mod_1318.get(0);
        mod_1351.put(0, t);
    endrule
    rule rule_1713;
        ChannelMessage t;
        t <- mod_1345.get(0);
        mod_1344.put(1, t);
    endrule
    rule rule_1714;
        ChannelMessage t;
        t <- mod_1350.get(0);
        mod_1320.put(1, t);
    endrule
    rule rule_1715;
        ChannelMessage t;
        t <- mod_1334.get(0);
        mod_1332.put(0, t);
    endrule
    rule rule_1716;
        ChannelMessage t;
        t <- mod_1321.get(0);
        mod_1322.put(0, t);
    endrule
    rule rule_1717;
        ChannelMessage t;
        t <- mod_1344.get(1);
        mod_1339.put(0, t);
    endrule
    rule rule_1718;
        ChannelMessage t;
        t <- mod_1313.get(0);
        mod_1314.put(0, t);
    endrule
    rule rule_1719;
        ChannelMessage t;
        t <- mod_1352.get(1);
        mod_1316.put(1, t);
    endrule
    rule rule_1720;
        ChannelMessage t;
        t <- mod_1346.get(1);
        mod_1321.put(1, t);
    endrule
    rule rule_1721;
        ChannelMessage t;
        t <- mod_1316.get(1);
        mod_1317.put(0, t);
    endrule
    rule rule_1722;
        ChannelMessage t;
        t <- mod_1326.get(0);
        mod_1327.put(0, t);
    endrule
    rule rule_1723;
        ChannelMessage t;
        t <- mod_1339.get(0);
        mod_1338.put(0, t);
    endrule
    rule rule_1724;
        ChannelMessage t;
        t <- mod_1315.get(0);
        mod_1316.put(0, t);
    endrule
    rule rule_1725;
        ChannelMessage t;
        t <- mod_1342.get(0);
        mod_1340.put(0, t);
    endrule
    rule rule_1726;
        ChannelMessage t;
        t <- mod_1335.get(0);
        mod_1334.put(0, t);
    endrule
    rule rule_1727;
        ChannelMessage t;
        t <- mod_1337.get(0);
        mod_1323.put(1, t);
    endrule
    rule rule_1728;
        ChannelMessage t;
        t <- mod_1319.get(1);
        mod_1320.put(0, t);
    endrule
    rule rule_1729;
        ChannelMessage t;
        t <- mod_1349.get(0);
        mod_1348.put(0, t);
    endrule
    rule rule_1730;
        ChannelMessage t;
        t <- mod_1351.get(0);
        mod_1318.put(1, t);
    endrule
    rule rule_1731;
        ChannelMessage t;
        t <- mod_1332.get(1);
        mod_1325.put(1, t);
    endrule
    rule rule_1732;
        ChannelMessage t;
        t <- mod_1325.get(0);
        mod_1326.put(0, t);
    endrule
    rule rule_1733;
        ChannelMessage t;
        t <- mod_1348.get(0);
        mod_1346.put(0, t);
    endrule
    rule rule_1734;
        ChannelMessage t;
        t <- mod_1352.get(0);
        mod_1352.put(1, t);
    endrule
    rule rule_1735;
        ChannelMessage t;
        t <- mod_1332.get(0);
        mod_1333.put(0, t);
    endrule
    rule rule_1736;
        ChannelMessage t;
        t <- mod_1320.get(1);
        mod_1321.put(0, t);
    endrule
    rule rule_1737;
        ChannelMessage t;
        t <- mod_1341.get(0);
        mod_1340.put(1, t);
    endrule
    rule rule_1738;
        ChannelMessage t;
        t <- mod_1328.get(0);
        mod_1330.put(0, t);
    endrule
    rule rule_1739;
        ChannelMessage t;
        t <- mod_1322.get(0);
        mod_1323.put(0, t);
    endrule
    rule rule_1740;
        ChannelMessage t;
        t <- mod_1331.get(0);
        mod_1331.put(1, t);
    endrule
    rule rule_1741;
        ChannelMessage t;
        t <- mod_1340.get(1);
        mod_1339.put(1, t);
    endrule
    rule rule_1742;
        ChannelMessage t;
        t <- mod_1319.get(0);
        mod_1344.put(0, t);
    endrule
    rule rule_1743;
        ChannelMessage t;
        t <- mod_1330.get(1);
        mod_1328.put(1, t);
    endrule
    rule rule_1744;
        ChannelMessage t;
        t <- mod_1316.get(0);
        mod_1352.put(0, t);
    endrule
    rule rule_1745;
        ChannelMessage t;
        t <- mod_1317.get(3);
        mod_1318.put(0, t);
    endrule
    rule rule_1746;
        ChannelMessage t;
        t <- mod_1314.get(0);
        mod_1315.put(0, t);
    endrule
    rule rule_1747;
        ChannelMessage t;
        t <- mod_1327.get(1);
        mod_1328.put(0, t);
    endrule
    rule rule_1748;
        ChannelMessage t;
        t <- mod_1343.get(0);
        mod_1342.put(0, t);
    endrule
    rule rule_1749;
        ChannelMessage t;
        t <- mod_1324.get(0);
        mod_1336.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1313.put(0, t);
        end
        if (i == 1) begin
            mod_1329.put(0, t);
        end
        if (i == 2) begin
            mod_1335.put(0, t);
        end
        if (i == 3) begin
            mod_1343.put(0, t);
        end
        if (i == 4) begin
            mod_1349.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_1317.get(0);
        end
        if (i == 2) begin
            t <- mod_1317.get(1);
        end
        if (i == 1) begin
            t <- mod_1317.get(2);
        end
        if (i == 3) begin
            t <- mod_1329.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6067 (Operation_IFC);
    Operation_IFC mod_1354_inner <- mkReshape(2, 64);
    Operation_IFC mod_1354 <- mkDebugOperation(mod_1354_inner, "mod_1354");
    Operation_IFC mod_1355_inner <- mkFlatten(1);
    Operation_IFC mod_1355 <- mkDebugOperation(mod_1355_inner, "mod_1355");
    Operation_IFC mod_1356_inner <- mkFlatten(2);
    Operation_IFC mod_1356 <- mkDebugOperation(mod_1356_inner, "mod_1356");
    Operation_IFC mod_1357_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1357 <- mkDebugOperation(mod_1357_inner, "mod_1357");
    Broadcast_IFC#(4) mod_1358_inner <- mkBroadcast(4);
    Operation_IFC mod_1358 <- mkDebugOperation(mod_1358_inner.op, "mod_1358");
    PMU_IFC mod_1359_bufferize <- mkPMU(2);
    Operation_IFC mod_1359_inner = mod_1359_bufferize.operation;
    Operation_IFC mod_1359 <- mkDebugOperation(mod_1359_inner, "mod_1359");
    Broadcast_IFC#(2) mod_1360_inner <- mkBroadcast(2);
    Operation_IFC mod_1360 <- mkDebugOperation(mod_1360_inner.op, "mod_1360");
    PMU_IFC mod_1361_bufferize <- mkPMU(1);
    Operation_IFC mod_1361_inner = mod_1361_bufferize.operation;
    Operation_IFC mod_1361 <- mkDebugOperation(mod_1361_inner, "mod_1361");
    Operation_IFC mod_1362_inner <- mkBinaryMap(1123, matmul_t_tile);
    Operation_IFC mod_1362 <- mkDebugOperation(mod_1362_inner, "mod_1362");
    Operation_IFC mod_1363_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1363 <- mkDebugOperation(mod_1363_inner, "mod_1363");
    Operation_IFC mod_1364_inner <- mkBinaryMap(1891, mul_tile);
    Operation_IFC mod_1364 <- mkDebugOperation(mod_1364_inner, "mod_1364");
    PMU_IFC mod_1365_bufferize <- mkPMU(1);
    Operation_IFC mod_1365_inner = mod_1365_bufferize.operation;
    Operation_IFC mod_1365 <- mkDebugOperation(mod_1365_inner, "mod_1365");
    Operation_IFC mod_1366_inner <- mkBinaryMap(2497, matmul_t_tile);
    Operation_IFC mod_1366 <- mkDebugOperation(mod_1366_inner, "mod_1366");
    Operation_IFC mod_1367_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1367 <- mkDebugOperation(mod_1367_inner, "mod_1367");
    Operation_IFC mod_1368_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1368 <- mkDebugOperation(mod_1368_inner, "mod_1368");
    Operation_IFC mod_1369_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1369 <- mkDebugOperation(mod_1369_inner, "mod_1369");
    Operation_IFC mod_1370_inner <- mkBinaryMap(2790, mul_tile);
    Operation_IFC mod_1370 <- mkDebugOperation(mod_1370_inner, "mod_1370");
    PMU_IFC mod_1371_bufferize <- mkPMU(1);
    Operation_IFC mod_1371_inner = mod_1371_bufferize.operation;
    Operation_IFC mod_1371 <- mkDebugOperation(mod_1371_inner, "mod_1371");
    PMU_IFC mod_1372_bufferize <- mkPMU(2);
    Operation_IFC mod_1372_inner = mod_1372_bufferize.operation;
    Operation_IFC mod_1372 <- mkDebugOperation(mod_1372_inner, "mod_1372");
    PMU_IFC mod_1373_bufferize <- mkPMU(2);
    Operation_IFC mod_1373_inner = mod_1373_bufferize.operation;
    Operation_IFC mod_1373 <- mkDebugOperation(mod_1373_inner, "mod_1373");
    Operation_IFC mod_1374_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1374 <- mkDebugOperation(mod_1374_inner, "mod_1374");
    Operation_IFC mod_1375_inner <- mkFlatten(1);
    Operation_IFC mod_1375 <- mkDebugOperation(mod_1375_inner, "mod_1375");
    Operation_IFC mod_1376_inner <- mkFlatten(0);
    Operation_IFC mod_1376 <- mkDebugOperation(mod_1376_inner, "mod_1376");
    Operation_IFC mod_1377_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1377 <- mkDebugOperation(mod_1377_inner, "mod_1377");
    Operation_IFC mod_1378_inner <- mkUnaryMap(1763, silu_tile);
    Operation_IFC mod_1378 <- mkDebugOperation(mod_1378_inner, "mod_1378");
    Operation_IFC mod_1379_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1379 <- mkDebugOperation(mod_1379_inner, "mod_1379");
    Operation_IFC mod_1380_inner <- mkBinaryMap(1635, matmul_t_tile);
    Operation_IFC mod_1380 <- mkDebugOperation(mod_1380_inner, "mod_1380");
    PMU_IFC mod_1381_bufferize <- mkPMU(2);
    Operation_IFC mod_1381_inner = mod_1381_bufferize.operation;
    Operation_IFC mod_1381 <- mkDebugOperation(mod_1381_inner, "mod_1381");
    Operation_IFC mod_1382_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1382 <- mkDebugOperation(mod_1382_inner, "mod_1382");
    Operation_IFC mod_1383_inner <- mkFlatten(1);
    Operation_IFC mod_1383 <- mkDebugOperation(mod_1383_inner, "mod_1383");
    Operation_IFC mod_1384_inner <- mkFlatten(0);
    Operation_IFC mod_1384 <- mkDebugOperation(mod_1384_inner, "mod_1384");
    PMU_IFC mod_1385_bufferize <- mkPMU(1);
    Operation_IFC mod_1385_inner = mod_1385_bufferize.operation;
    Operation_IFC mod_1385 <- mkDebugOperation(mod_1385_inner, "mod_1385");
    Operation_IFC mod_1386_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1386 <- mkDebugOperation(mod_1386_inner, "mod_1386");
    PMU_IFC mod_1387_bufferize <- mkPMU(2);
    Operation_IFC mod_1387_inner = mod_1387_bufferize.operation;
    Operation_IFC mod_1387 <- mkDebugOperation(mod_1387_inner, "mod_1387");
    Operation_IFC mod_1388_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1388 <- mkDebugOperation(mod_1388_inner, "mod_1388");
    Operation_IFC mod_1389_inner <- mkFlatten(1);
    Operation_IFC mod_1389 <- mkDebugOperation(mod_1389_inner, "mod_1389");
    Operation_IFC mod_1390_inner <- mkFlatten(0);
    Operation_IFC mod_1390 <- mkDebugOperation(mod_1390_inner, "mod_1390");
    Operation_IFC mod_1391_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1391 <- mkDebugOperation(mod_1391_inner, "mod_1391");
    Operation_IFC mod_1392_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1392 <- mkDebugOperation(mod_1392_inner, "mod_1392");
    PMU_IFC mod_1393_bufferize <- mkPMU(2);
    Operation_IFC mod_1393_inner = mod_1393_bufferize.operation;
    Operation_IFC mod_1393 <- mkDebugOperation(mod_1393_inner, "mod_1393");
    rule rule_1750;
        ChannelMessage t;
        t <- mod_1387.get(1);
        mod_1362.put(1, t);
    endrule
    rule rule_1751;
        ChannelMessage t;
        t <- mod_1369.get(1);
        mod_1370.put(1, t);
    endrule
    rule rule_1752;
        ChannelMessage t;
        t <- mod_1373.get(1);
        mod_1366.put(1, t);
    endrule
    rule rule_1753;
        ChannelMessage t;
        t <- mod_1374.get(0);
        mod_1373.put(1, t);
    endrule
    rule rule_1754;
        ChannelMessage t;
        t <- mod_1391.get(0);
        mod_1361.put(1, t);
    endrule
    rule rule_1755;
        ChannelMessage t;
        t <- mod_1373.get(0);
        mod_1374.put(0, t);
    endrule
    rule rule_1756;
        ChannelMessage t;
        t <- mod_1354.get(0);
        mod_1355.put(0, t);
    endrule
    rule rule_1757;
        ChannelMessage t;
        t <- mod_1372.get(1);
        mod_1368.put(1, t);
    endrule
    rule rule_1758;
        ChannelMessage t;
        t <- mod_1361.get(1);
        mod_1362.put(0, t);
    endrule
    rule rule_1759;
        ChannelMessage t;
        t <- mod_1365.get(0);
        mod_1377.put(0, t);
    endrule
    rule rule_1760;
        ChannelMessage t;
        t <- mod_1377.get(0);
        mod_1365.put(1, t);
    endrule
    rule rule_1761;
        ChannelMessage t;
        t <- mod_1369.get(0);
        mod_1371.put(0, t);
    endrule
    rule rule_1762;
        ChannelMessage t;
        t <- mod_1359.get(1);
        mod_1360.put(0, t);
    endrule
    rule rule_1763;
        ChannelMessage t;
        t <- mod_1363.get(0);
        mod_1364.put(0, t);
    endrule
    rule rule_1764;
        ChannelMessage t;
        t <- mod_1364.get(0);
        mod_1365.put(0, t);
    endrule
    rule rule_1765;
        ChannelMessage t;
        t <- mod_1371.get(1);
        mod_1369.put(1, t);
    endrule
    rule rule_1766;
        ChannelMessage t;
        t <- mod_1375.get(0);
        mod_1373.put(0, t);
    endrule
    rule rule_1767;
        ChannelMessage t;
        t <- mod_1356.get(0);
        mod_1357.put(0, t);
    endrule
    rule rule_1768;
        ChannelMessage t;
        t <- mod_1382.get(0);
        mod_1381.put(1, t);
    endrule
    rule rule_1769;
        ChannelMessage t;
        t <- mod_1392.get(0);
        mod_1359.put(1, t);
    endrule
    rule rule_1770;
        ChannelMessage t;
        t <- mod_1371.get(0);
        mod_1371.put(1, t);
    endrule
    rule rule_1771;
        ChannelMessage t;
        t <- mod_1387.get(0);
        mod_1388.put(0, t);
    endrule
    rule rule_1772;
        ChannelMessage t;
        t <- mod_1379.get(0);
        mod_1378.put(0, t);
    endrule
    rule rule_1773;
        ChannelMessage t;
        t <- mod_1384.get(0);
        mod_1383.put(0, t);
    endrule
    rule rule_1774;
        ChannelMessage t;
        t <- mod_1378.get(0);
        mod_1364.put(1, t);
    endrule
    rule rule_1775;
        ChannelMessage t;
        t <- mod_1372.get(0);
        mod_1372.put(1, t);
    endrule
    rule rule_1776;
        ChannelMessage t;
        t <- mod_1368.get(1);
        mod_1369.put(0, t);
    endrule
    rule rule_1777;
        ChannelMessage t;
        t <- mod_1360.get(0);
        mod_1385.put(0, t);
    endrule
    rule rule_1778;
        ChannelMessage t;
        t <- mod_1381.get(0);
        mod_1382.put(0, t);
    endrule
    rule rule_1779;
        ChannelMessage t;
        t <- mod_1393.get(1);
        mod_1357.put(1, t);
    endrule
    rule rule_1780;
        ChannelMessage t;
        t <- mod_1388.get(0);
        mod_1387.put(1, t);
    endrule
    rule rule_1781;
        ChannelMessage t;
        t <- mod_1385.get(0);
        mod_1386.put(0, t);
    endrule
    rule rule_1782;
        ChannelMessage t;
        t <- mod_1357.get(1);
        mod_1358.put(0, t);
    endrule
    rule rule_1783;
        ChannelMessage t;
        t <- mod_1380.get(0);
        mod_1379.put(0, t);
    endrule
    rule rule_1784;
        ChannelMessage t;
        t <- mod_1389.get(0);
        mod_1387.put(0, t);
    endrule
    rule rule_1785;
        ChannelMessage t;
        t <- mod_1390.get(0);
        mod_1389.put(0, t);
    endrule
    rule rule_1786;
        ChannelMessage t;
        t <- mod_1393.get(0);
        mod_1393.put(1, t);
    endrule
    rule rule_1787;
        ChannelMessage t;
        t <- mod_1359.get(0);
        mod_1392.put(0, t);
    endrule
    rule rule_1788;
        ChannelMessage t;
        t <- mod_1360.get(1);
        mod_1361.put(0, t);
    endrule
    rule rule_1789;
        ChannelMessage t;
        t <- mod_1358.get(3);
        mod_1359.put(0, t);
    endrule
    rule rule_1790;
        ChannelMessage t;
        t <- mod_1366.get(0);
        mod_1367.put(0, t);
    endrule
    rule rule_1791;
        ChannelMessage t;
        t <- mod_1381.get(1);
        mod_1380.put(1, t);
    endrule
    rule rule_1792;
        ChannelMessage t;
        t <- mod_1386.get(0);
        mod_1385.put(1, t);
    endrule
    rule rule_1793;
        ChannelMessage t;
        t <- mod_1367.get(0);
        mod_1368.put(0, t);
    endrule
    rule rule_1794;
        ChannelMessage t;
        t <- mod_1361.get(0);
        mod_1391.put(0, t);
    endrule
    rule rule_1795;
        ChannelMessage t;
        t <- mod_1357.get(0);
        mod_1393.put(0, t);
    endrule
    rule rule_1796;
        ChannelMessage t;
        t <- mod_1383.get(0);
        mod_1381.put(0, t);
    endrule
    rule rule_1797;
        ChannelMessage t;
        t <- mod_1385.get(1);
        mod_1380.put(0, t);
    endrule
    rule rule_1798;
        ChannelMessage t;
        t <- mod_1365.get(1);
        mod_1366.put(0, t);
    endrule
    rule rule_1799;
        ChannelMessage t;
        t <- mod_1376.get(0);
        mod_1375.put(0, t);
    endrule
    rule rule_1800;
        ChannelMessage t;
        t <- mod_1355.get(0);
        mod_1356.put(0, t);
    endrule
    rule rule_1801;
        ChannelMessage t;
        t <- mod_1362.get(0);
        mod_1363.put(0, t);
    endrule
    rule rule_1802;
        ChannelMessage t;
        t <- mod_1368.get(0);
        mod_1372.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1354.put(0, t);
        end
        if (i == 1) begin
            mod_1370.put(0, t);
        end
        if (i == 2) begin
            mod_1376.put(0, t);
        end
        if (i == 3) begin
            mod_1384.put(0, t);
        end
        if (i == 4) begin
            mod_1390.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 2) begin
            t <- mod_1358.get(0);
        end
        if (i == 3) begin
            t <- mod_1358.get(1);
        end
        if (i == 1) begin
            t <- mod_1358.get(2);
        end
        if (i == 0) begin
            t <- mod_1370.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6068 (Operation_IFC);
    Operation_IFC mod_1395_inner <- mkReshape(2, 64);
    Operation_IFC mod_1395 <- mkDebugOperation(mod_1395_inner, "mod_1395");
    Operation_IFC mod_1396_inner <- mkFlatten(1);
    Operation_IFC mod_1396 <- mkDebugOperation(mod_1396_inner, "mod_1396");
    Operation_IFC mod_1397_inner <- mkFlatten(2);
    Operation_IFC mod_1397 <- mkDebugOperation(mod_1397_inner, "mod_1397");
    Operation_IFC mod_1398_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1398 <- mkDebugOperation(mod_1398_inner, "mod_1398");
    Broadcast_IFC#(4) mod_1399_inner <- mkBroadcast(4);
    Operation_IFC mod_1399 <- mkDebugOperation(mod_1399_inner.op, "mod_1399");
    PMU_IFC mod_1400_bufferize <- mkPMU(2);
    Operation_IFC mod_1400_inner = mod_1400_bufferize.operation;
    Operation_IFC mod_1400 <- mkDebugOperation(mod_1400_inner, "mod_1400");
    Broadcast_IFC#(2) mod_1401_inner <- mkBroadcast(2);
    Operation_IFC mod_1401 <- mkDebugOperation(mod_1401_inner.op, "mod_1401");
    PMU_IFC mod_1402_bufferize <- mkPMU(1);
    Operation_IFC mod_1402_inner = mod_1402_bufferize.operation;
    Operation_IFC mod_1402 <- mkDebugOperation(mod_1402_inner, "mod_1402");
    Operation_IFC mod_1403_inner <- mkBinaryMap(1122, matmul_t_tile);
    Operation_IFC mod_1403 <- mkDebugOperation(mod_1403_inner, "mod_1403");
    Operation_IFC mod_1404_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1404 <- mkDebugOperation(mod_1404_inner, "mod_1404");
    Operation_IFC mod_1405_inner <- mkBinaryMap(1890, mul_tile);
    Operation_IFC mod_1405 <- mkDebugOperation(mod_1405_inner, "mod_1405");
    PMU_IFC mod_1406_bufferize <- mkPMU(1);
    Operation_IFC mod_1406_inner = mod_1406_bufferize.operation;
    Operation_IFC mod_1406 <- mkDebugOperation(mod_1406_inner, "mod_1406");
    Operation_IFC mod_1407_inner <- mkBinaryMap(2495, matmul_t_tile);
    Operation_IFC mod_1407 <- mkDebugOperation(mod_1407_inner, "mod_1407");
    Operation_IFC mod_1408_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1408 <- mkDebugOperation(mod_1408_inner, "mod_1408");
    Operation_IFC mod_1409_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1409 <- mkDebugOperation(mod_1409_inner, "mod_1409");
    Operation_IFC mod_1410_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1410 <- mkDebugOperation(mod_1410_inner, "mod_1410");
    Operation_IFC mod_1411_inner <- mkBinaryMap(2789, mul_tile);
    Operation_IFC mod_1411 <- mkDebugOperation(mod_1411_inner, "mod_1411");
    PMU_IFC mod_1412_bufferize <- mkPMU(1);
    Operation_IFC mod_1412_inner = mod_1412_bufferize.operation;
    Operation_IFC mod_1412 <- mkDebugOperation(mod_1412_inner, "mod_1412");
    PMU_IFC mod_1413_bufferize <- mkPMU(2);
    Operation_IFC mod_1413_inner = mod_1413_bufferize.operation;
    Operation_IFC mod_1413 <- mkDebugOperation(mod_1413_inner, "mod_1413");
    PMU_IFC mod_1414_bufferize <- mkPMU(2);
    Operation_IFC mod_1414_inner = mod_1414_bufferize.operation;
    Operation_IFC mod_1414 <- mkDebugOperation(mod_1414_inner, "mod_1414");
    Operation_IFC mod_1415_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1415 <- mkDebugOperation(mod_1415_inner, "mod_1415");
    Operation_IFC mod_1416_inner <- mkFlatten(1);
    Operation_IFC mod_1416 <- mkDebugOperation(mod_1416_inner, "mod_1416");
    Operation_IFC mod_1417_inner <- mkFlatten(0);
    Operation_IFC mod_1417 <- mkDebugOperation(mod_1417_inner, "mod_1417");
    Operation_IFC mod_1418_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1418 <- mkDebugOperation(mod_1418_inner, "mod_1418");
    Operation_IFC mod_1419_inner <- mkUnaryMap(1762, silu_tile);
    Operation_IFC mod_1419 <- mkDebugOperation(mod_1419_inner, "mod_1419");
    Operation_IFC mod_1420_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1420 <- mkDebugOperation(mod_1420_inner, "mod_1420");
    Operation_IFC mod_1421_inner <- mkBinaryMap(1634, matmul_t_tile);
    Operation_IFC mod_1421 <- mkDebugOperation(mod_1421_inner, "mod_1421");
    PMU_IFC mod_1422_bufferize <- mkPMU(2);
    Operation_IFC mod_1422_inner = mod_1422_bufferize.operation;
    Operation_IFC mod_1422 <- mkDebugOperation(mod_1422_inner, "mod_1422");
    Operation_IFC mod_1423_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1423 <- mkDebugOperation(mod_1423_inner, "mod_1423");
    Operation_IFC mod_1424_inner <- mkFlatten(1);
    Operation_IFC mod_1424 <- mkDebugOperation(mod_1424_inner, "mod_1424");
    Operation_IFC mod_1425_inner <- mkFlatten(0);
    Operation_IFC mod_1425 <- mkDebugOperation(mod_1425_inner, "mod_1425");
    PMU_IFC mod_1426_bufferize <- mkPMU(1);
    Operation_IFC mod_1426_inner = mod_1426_bufferize.operation;
    Operation_IFC mod_1426 <- mkDebugOperation(mod_1426_inner, "mod_1426");
    Operation_IFC mod_1427_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1427 <- mkDebugOperation(mod_1427_inner, "mod_1427");
    PMU_IFC mod_1428_bufferize <- mkPMU(2);
    Operation_IFC mod_1428_inner = mod_1428_bufferize.operation;
    Operation_IFC mod_1428 <- mkDebugOperation(mod_1428_inner, "mod_1428");
    Operation_IFC mod_1429_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1429 <- mkDebugOperation(mod_1429_inner, "mod_1429");
    Operation_IFC mod_1430_inner <- mkFlatten(1);
    Operation_IFC mod_1430 <- mkDebugOperation(mod_1430_inner, "mod_1430");
    Operation_IFC mod_1431_inner <- mkFlatten(0);
    Operation_IFC mod_1431 <- mkDebugOperation(mod_1431_inner, "mod_1431");
    Operation_IFC mod_1432_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1432 <- mkDebugOperation(mod_1432_inner, "mod_1432");
    Operation_IFC mod_1433_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1433 <- mkDebugOperation(mod_1433_inner, "mod_1433");
    PMU_IFC mod_1434_bufferize <- mkPMU(2);
    Operation_IFC mod_1434_inner = mod_1434_bufferize.operation;
    Operation_IFC mod_1434 <- mkDebugOperation(mod_1434_inner, "mod_1434");
    rule rule_1803;
        ChannelMessage t;
        t <- mod_1432.get(0);
        mod_1402.put(1, t);
    endrule
    rule rule_1804;
        ChannelMessage t;
        t <- mod_1414.get(1);
        mod_1407.put(1, t);
    endrule
    rule rule_1805;
        ChannelMessage t;
        t <- mod_1400.get(0);
        mod_1433.put(0, t);
    endrule
    rule rule_1806;
        ChannelMessage t;
        t <- mod_1405.get(0);
        mod_1406.put(0, t);
    endrule
    rule rule_1807;
        ChannelMessage t;
        t <- mod_1433.get(0);
        mod_1400.put(1, t);
    endrule
    rule rule_1808;
        ChannelMessage t;
        t <- mod_1434.get(1);
        mod_1398.put(1, t);
    endrule
    rule rule_1809;
        ChannelMessage t;
        t <- mod_1399.get(3);
        mod_1400.put(0, t);
    endrule
    rule rule_1810;
        ChannelMessage t;
        t <- mod_1407.get(0);
        mod_1408.put(0, t);
    endrule
    rule rule_1811;
        ChannelMessage t;
        t <- mod_1406.get(0);
        mod_1418.put(0, t);
    endrule
    rule rule_1812;
        ChannelMessage t;
        t <- mod_1412.get(1);
        mod_1410.put(1, t);
    endrule
    rule rule_1813;
        ChannelMessage t;
        t <- mod_1404.get(0);
        mod_1405.put(0, t);
    endrule
    rule rule_1814;
        ChannelMessage t;
        t <- mod_1429.get(0);
        mod_1428.put(1, t);
    endrule
    rule rule_1815;
        ChannelMessage t;
        t <- mod_1408.get(0);
        mod_1409.put(0, t);
    endrule
    rule rule_1816;
        ChannelMessage t;
        t <- mod_1409.get(0);
        mod_1413.put(0, t);
    endrule
    rule rule_1817;
        ChannelMessage t;
        t <- mod_1401.get(1);
        mod_1402.put(0, t);
    endrule
    rule rule_1818;
        ChannelMessage t;
        t <- mod_1397.get(0);
        mod_1398.put(0, t);
    endrule
    rule rule_1819;
        ChannelMessage t;
        t <- mod_1396.get(0);
        mod_1397.put(0, t);
    endrule
    rule rule_1820;
        ChannelMessage t;
        t <- mod_1395.get(0);
        mod_1396.put(0, t);
    endrule
    rule rule_1821;
        ChannelMessage t;
        t <- mod_1410.get(1);
        mod_1411.put(1, t);
    endrule
    rule rule_1822;
        ChannelMessage t;
        t <- mod_1423.get(0);
        mod_1422.put(1, t);
    endrule
    rule rule_1823;
        ChannelMessage t;
        t <- mod_1426.get(1);
        mod_1421.put(0, t);
    endrule
    rule rule_1824;
        ChannelMessage t;
        t <- mod_1403.get(0);
        mod_1404.put(0, t);
    endrule
    rule rule_1825;
        ChannelMessage t;
        t <- mod_1422.get(1);
        mod_1421.put(1, t);
    endrule
    rule rule_1826;
        ChannelMessage t;
        t <- mod_1428.get(1);
        mod_1403.put(1, t);
    endrule
    rule rule_1827;
        ChannelMessage t;
        t <- mod_1421.get(0);
        mod_1420.put(0, t);
    endrule
    rule rule_1828;
        ChannelMessage t;
        t <- mod_1414.get(0);
        mod_1415.put(0, t);
    endrule
    rule rule_1829;
        ChannelMessage t;
        t <- mod_1420.get(0);
        mod_1419.put(0, t);
    endrule
    rule rule_1830;
        ChannelMessage t;
        t <- mod_1410.get(0);
        mod_1412.put(0, t);
    endrule
    rule rule_1831;
        ChannelMessage t;
        t <- mod_1413.get(0);
        mod_1413.put(1, t);
    endrule
    rule rule_1832;
        ChannelMessage t;
        t <- mod_1400.get(1);
        mod_1401.put(0, t);
    endrule
    rule rule_1833;
        ChannelMessage t;
        t <- mod_1398.get(1);
        mod_1399.put(0, t);
    endrule
    rule rule_1834;
        ChannelMessage t;
        t <- mod_1418.get(0);
        mod_1406.put(1, t);
    endrule
    rule rule_1835;
        ChannelMessage t;
        t <- mod_1398.get(0);
        mod_1434.put(0, t);
    endrule
    rule rule_1836;
        ChannelMessage t;
        t <- mod_1426.get(0);
        mod_1427.put(0, t);
    endrule
    rule rule_1837;
        ChannelMessage t;
        t <- mod_1415.get(0);
        mod_1414.put(1, t);
    endrule
    rule rule_1838;
        ChannelMessage t;
        t <- mod_1402.get(0);
        mod_1432.put(0, t);
    endrule
    rule rule_1839;
        ChannelMessage t;
        t <- mod_1402.get(1);
        mod_1403.put(0, t);
    endrule
    rule rule_1840;
        ChannelMessage t;
        t <- mod_1427.get(0);
        mod_1426.put(1, t);
    endrule
    rule rule_1841;
        ChannelMessage t;
        t <- mod_1428.get(0);
        mod_1429.put(0, t);
    endrule
    rule rule_1842;
        ChannelMessage t;
        t <- mod_1406.get(1);
        mod_1407.put(0, t);
    endrule
    rule rule_1843;
        ChannelMessage t;
        t <- mod_1413.get(1);
        mod_1409.put(1, t);
    endrule
    rule rule_1844;
        ChannelMessage t;
        t <- mod_1430.get(0);
        mod_1428.put(0, t);
    endrule
    rule rule_1845;
        ChannelMessage t;
        t <- mod_1422.get(0);
        mod_1423.put(0, t);
    endrule
    rule rule_1846;
        ChannelMessage t;
        t <- mod_1401.get(0);
        mod_1426.put(0, t);
    endrule
    rule rule_1847;
        ChannelMessage t;
        t <- mod_1409.get(1);
        mod_1410.put(0, t);
    endrule
    rule rule_1848;
        ChannelMessage t;
        t <- mod_1424.get(0);
        mod_1422.put(0, t);
    endrule
    rule rule_1849;
        ChannelMessage t;
        t <- mod_1416.get(0);
        mod_1414.put(0, t);
    endrule
    rule rule_1850;
        ChannelMessage t;
        t <- mod_1431.get(0);
        mod_1430.put(0, t);
    endrule
    rule rule_1851;
        ChannelMessage t;
        t <- mod_1425.get(0);
        mod_1424.put(0, t);
    endrule
    rule rule_1852;
        ChannelMessage t;
        t <- mod_1419.get(0);
        mod_1405.put(1, t);
    endrule
    rule rule_1853;
        ChannelMessage t;
        t <- mod_1412.get(0);
        mod_1412.put(1, t);
    endrule
    rule rule_1854;
        ChannelMessage t;
        t <- mod_1434.get(0);
        mod_1434.put(1, t);
    endrule
    rule rule_1855;
        ChannelMessage t;
        t <- mod_1417.get(0);
        mod_1416.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1395.put(0, t);
        end
        if (i == 1) begin
            mod_1411.put(0, t);
        end
        if (i == 2) begin
            mod_1417.put(0, t);
        end
        if (i == 3) begin
            mod_1425.put(0, t);
        end
        if (i == 4) begin
            mod_1431.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_1399.get(0);
        end
        if (i == 0) begin
            t <- mod_1399.get(1);
        end
        if (i == 1) begin
            t <- mod_1399.get(2);
        end
        if (i == 2) begin
            t <- mod_1411.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6069 (Operation_IFC);
    Operation_IFC mod_1436_inner <- mkReshape(2, 64);
    Operation_IFC mod_1436 <- mkDebugOperation(mod_1436_inner, "mod_1436");
    Operation_IFC mod_1437_inner <- mkFlatten(1);
    Operation_IFC mod_1437 <- mkDebugOperation(mod_1437_inner, "mod_1437");
    Operation_IFC mod_1438_inner <- mkFlatten(2);
    Operation_IFC mod_1438 <- mkDebugOperation(mod_1438_inner, "mod_1438");
    Operation_IFC mod_1439_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1439 <- mkDebugOperation(mod_1439_inner, "mod_1439");
    Broadcast_IFC#(4) mod_1440_inner <- mkBroadcast(4);
    Operation_IFC mod_1440 <- mkDebugOperation(mod_1440_inner.op, "mod_1440");
    PMU_IFC mod_1441_bufferize <- mkPMU(2);
    Operation_IFC mod_1441_inner = mod_1441_bufferize.operation;
    Operation_IFC mod_1441 <- mkDebugOperation(mod_1441_inner, "mod_1441");
    Broadcast_IFC#(2) mod_1442_inner <- mkBroadcast(2);
    Operation_IFC mod_1442 <- mkDebugOperation(mod_1442_inner.op, "mod_1442");
    PMU_IFC mod_1443_bufferize <- mkPMU(1);
    Operation_IFC mod_1443_inner = mod_1443_bufferize.operation;
    Operation_IFC mod_1443 <- mkDebugOperation(mod_1443_inner, "mod_1443");
    Operation_IFC mod_1444_inner <- mkBinaryMap(1121, matmul_t_tile);
    Operation_IFC mod_1444 <- mkDebugOperation(mod_1444_inner, "mod_1444");
    Operation_IFC mod_1445_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1445 <- mkDebugOperation(mod_1445_inner, "mod_1445");
    Operation_IFC mod_1446_inner <- mkBinaryMap(1889, mul_tile);
    Operation_IFC mod_1446 <- mkDebugOperation(mod_1446_inner, "mod_1446");
    PMU_IFC mod_1447_bufferize <- mkPMU(1);
    Operation_IFC mod_1447_inner = mod_1447_bufferize.operation;
    Operation_IFC mod_1447 <- mkDebugOperation(mod_1447_inner, "mod_1447");
    Operation_IFC mod_1448_inner <- mkBinaryMap(2493, matmul_t_tile);
    Operation_IFC mod_1448 <- mkDebugOperation(mod_1448_inner, "mod_1448");
    Operation_IFC mod_1449_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1449 <- mkDebugOperation(mod_1449_inner, "mod_1449");
    Operation_IFC mod_1450_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1450 <- mkDebugOperation(mod_1450_inner, "mod_1450");
    Operation_IFC mod_1451_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1451 <- mkDebugOperation(mod_1451_inner, "mod_1451");
    Operation_IFC mod_1452_inner <- mkBinaryMap(2788, mul_tile);
    Operation_IFC mod_1452 <- mkDebugOperation(mod_1452_inner, "mod_1452");
    PMU_IFC mod_1453_bufferize <- mkPMU(1);
    Operation_IFC mod_1453_inner = mod_1453_bufferize.operation;
    Operation_IFC mod_1453 <- mkDebugOperation(mod_1453_inner, "mod_1453");
    PMU_IFC mod_1454_bufferize <- mkPMU(2);
    Operation_IFC mod_1454_inner = mod_1454_bufferize.operation;
    Operation_IFC mod_1454 <- mkDebugOperation(mod_1454_inner, "mod_1454");
    PMU_IFC mod_1455_bufferize <- mkPMU(2);
    Operation_IFC mod_1455_inner = mod_1455_bufferize.operation;
    Operation_IFC mod_1455 <- mkDebugOperation(mod_1455_inner, "mod_1455");
    Operation_IFC mod_1456_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1456 <- mkDebugOperation(mod_1456_inner, "mod_1456");
    Operation_IFC mod_1457_inner <- mkFlatten(1);
    Operation_IFC mod_1457 <- mkDebugOperation(mod_1457_inner, "mod_1457");
    Operation_IFC mod_1458_inner <- mkFlatten(0);
    Operation_IFC mod_1458 <- mkDebugOperation(mod_1458_inner, "mod_1458");
    Operation_IFC mod_1459_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1459 <- mkDebugOperation(mod_1459_inner, "mod_1459");
    Operation_IFC mod_1460_inner <- mkUnaryMap(1761, silu_tile);
    Operation_IFC mod_1460 <- mkDebugOperation(mod_1460_inner, "mod_1460");
    Operation_IFC mod_1461_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1461 <- mkDebugOperation(mod_1461_inner, "mod_1461");
    Operation_IFC mod_1462_inner <- mkBinaryMap(1633, matmul_t_tile);
    Operation_IFC mod_1462 <- mkDebugOperation(mod_1462_inner, "mod_1462");
    PMU_IFC mod_1463_bufferize <- mkPMU(2);
    Operation_IFC mod_1463_inner = mod_1463_bufferize.operation;
    Operation_IFC mod_1463 <- mkDebugOperation(mod_1463_inner, "mod_1463");
    Operation_IFC mod_1464_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1464 <- mkDebugOperation(mod_1464_inner, "mod_1464");
    Operation_IFC mod_1465_inner <- mkFlatten(1);
    Operation_IFC mod_1465 <- mkDebugOperation(mod_1465_inner, "mod_1465");
    Operation_IFC mod_1466_inner <- mkFlatten(0);
    Operation_IFC mod_1466 <- mkDebugOperation(mod_1466_inner, "mod_1466");
    PMU_IFC mod_1467_bufferize <- mkPMU(1);
    Operation_IFC mod_1467_inner = mod_1467_bufferize.operation;
    Operation_IFC mod_1467 <- mkDebugOperation(mod_1467_inner, "mod_1467");
    Operation_IFC mod_1468_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1468 <- mkDebugOperation(mod_1468_inner, "mod_1468");
    PMU_IFC mod_1469_bufferize <- mkPMU(2);
    Operation_IFC mod_1469_inner = mod_1469_bufferize.operation;
    Operation_IFC mod_1469 <- mkDebugOperation(mod_1469_inner, "mod_1469");
    Operation_IFC mod_1470_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1470 <- mkDebugOperation(mod_1470_inner, "mod_1470");
    Operation_IFC mod_1471_inner <- mkFlatten(1);
    Operation_IFC mod_1471 <- mkDebugOperation(mod_1471_inner, "mod_1471");
    Operation_IFC mod_1472_inner <- mkFlatten(0);
    Operation_IFC mod_1472 <- mkDebugOperation(mod_1472_inner, "mod_1472");
    Operation_IFC mod_1473_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1473 <- mkDebugOperation(mod_1473_inner, "mod_1473");
    Operation_IFC mod_1474_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1474 <- mkDebugOperation(mod_1474_inner, "mod_1474");
    PMU_IFC mod_1475_bufferize <- mkPMU(2);
    Operation_IFC mod_1475_inner = mod_1475_bufferize.operation;
    Operation_IFC mod_1475 <- mkDebugOperation(mod_1475_inner, "mod_1475");
    rule rule_1856;
        ChannelMessage t;
        t <- mod_1474.get(0);
        mod_1441.put(1, t);
    endrule
    rule rule_1857;
        ChannelMessage t;
        t <- mod_1440.get(3);
        mod_1441.put(0, t);
    endrule
    rule rule_1858;
        ChannelMessage t;
        t <- mod_1454.get(0);
        mod_1454.put(1, t);
    endrule
    rule rule_1859;
        ChannelMessage t;
        t <- mod_1449.get(0);
        mod_1450.put(0, t);
    endrule
    rule rule_1860;
        ChannelMessage t;
        t <- mod_1463.get(0);
        mod_1464.put(0, t);
    endrule
    rule rule_1861;
        ChannelMessage t;
        t <- mod_1463.get(1);
        mod_1462.put(1, t);
    endrule
    rule rule_1862;
        ChannelMessage t;
        t <- mod_1455.get(0);
        mod_1456.put(0, t);
    endrule
    rule rule_1863;
        ChannelMessage t;
        t <- mod_1447.get(0);
        mod_1459.put(0, t);
    endrule
    rule rule_1864;
        ChannelMessage t;
        t <- mod_1461.get(0);
        mod_1460.put(0, t);
    endrule
    rule rule_1865;
        ChannelMessage t;
        t <- mod_1453.get(0);
        mod_1453.put(1, t);
    endrule
    rule rule_1866;
        ChannelMessage t;
        t <- mod_1438.get(0);
        mod_1439.put(0, t);
    endrule
    rule rule_1867;
        ChannelMessage t;
        t <- mod_1445.get(0);
        mod_1446.put(0, t);
    endrule
    rule rule_1868;
        ChannelMessage t;
        t <- mod_1441.get(0);
        mod_1474.put(0, t);
    endrule
    rule rule_1869;
        ChannelMessage t;
        t <- mod_1472.get(0);
        mod_1471.put(0, t);
    endrule
    rule rule_1870;
        ChannelMessage t;
        t <- mod_1450.get(0);
        mod_1454.put(0, t);
    endrule
    rule rule_1871;
        ChannelMessage t;
        t <- mod_1467.get(0);
        mod_1468.put(0, t);
    endrule
    rule rule_1872;
        ChannelMessage t;
        t <- mod_1475.get(1);
        mod_1439.put(1, t);
    endrule
    rule rule_1873;
        ChannelMessage t;
        t <- mod_1451.get(1);
        mod_1452.put(1, t);
    endrule
    rule rule_1874;
        ChannelMessage t;
        t <- mod_1460.get(0);
        mod_1446.put(1, t);
    endrule
    rule rule_1875;
        ChannelMessage t;
        t <- mod_1442.get(0);
        mod_1467.put(0, t);
    endrule
    rule rule_1876;
        ChannelMessage t;
        t <- mod_1457.get(0);
        mod_1455.put(0, t);
    endrule
    rule rule_1877;
        ChannelMessage t;
        t <- mod_1473.get(0);
        mod_1443.put(1, t);
    endrule
    rule rule_1878;
        ChannelMessage t;
        t <- mod_1439.get(1);
        mod_1440.put(0, t);
    endrule
    rule rule_1879;
        ChannelMessage t;
        t <- mod_1455.get(1);
        mod_1448.put(1, t);
    endrule
    rule rule_1880;
        ChannelMessage t;
        t <- mod_1442.get(1);
        mod_1443.put(0, t);
    endrule
    rule rule_1881;
        ChannelMessage t;
        t <- mod_1446.get(0);
        mod_1447.put(0, t);
    endrule
    rule rule_1882;
        ChannelMessage t;
        t <- mod_1441.get(1);
        mod_1442.put(0, t);
    endrule
    rule rule_1883;
        ChannelMessage t;
        t <- mod_1450.get(1);
        mod_1451.put(0, t);
    endrule
    rule rule_1884;
        ChannelMessage t;
        t <- mod_1443.get(0);
        mod_1473.put(0, t);
    endrule
    rule rule_1885;
        ChannelMessage t;
        t <- mod_1470.get(0);
        mod_1469.put(1, t);
    endrule
    rule rule_1886;
        ChannelMessage t;
        t <- mod_1465.get(0);
        mod_1463.put(0, t);
    endrule
    rule rule_1887;
        ChannelMessage t;
        t <- mod_1462.get(0);
        mod_1461.put(0, t);
    endrule
    rule rule_1888;
        ChannelMessage t;
        t <- mod_1475.get(0);
        mod_1475.put(1, t);
    endrule
    rule rule_1889;
        ChannelMessage t;
        t <- mod_1471.get(0);
        mod_1469.put(0, t);
    endrule
    rule rule_1890;
        ChannelMessage t;
        t <- mod_1436.get(0);
        mod_1437.put(0, t);
    endrule
    rule rule_1891;
        ChannelMessage t;
        t <- mod_1437.get(0);
        mod_1438.put(0, t);
    endrule
    rule rule_1892;
        ChannelMessage t;
        t <- mod_1444.get(0);
        mod_1445.put(0, t);
    endrule
    rule rule_1893;
        ChannelMessage t;
        t <- mod_1448.get(0);
        mod_1449.put(0, t);
    endrule
    rule rule_1894;
        ChannelMessage t;
        t <- mod_1453.get(1);
        mod_1451.put(1, t);
    endrule
    rule rule_1895;
        ChannelMessage t;
        t <- mod_1451.get(0);
        mod_1453.put(0, t);
    endrule
    rule rule_1896;
        ChannelMessage t;
        t <- mod_1458.get(0);
        mod_1457.put(0, t);
    endrule
    rule rule_1897;
        ChannelMessage t;
        t <- mod_1459.get(0);
        mod_1447.put(1, t);
    endrule
    rule rule_1898;
        ChannelMessage t;
        t <- mod_1464.get(0);
        mod_1463.put(1, t);
    endrule
    rule rule_1899;
        ChannelMessage t;
        t <- mod_1443.get(1);
        mod_1444.put(0, t);
    endrule
    rule rule_1900;
        ChannelMessage t;
        t <- mod_1468.get(0);
        mod_1467.put(1, t);
    endrule
    rule rule_1901;
        ChannelMessage t;
        t <- mod_1467.get(1);
        mod_1462.put(0, t);
    endrule
    rule rule_1902;
        ChannelMessage t;
        t <- mod_1454.get(1);
        mod_1450.put(1, t);
    endrule
    rule rule_1903;
        ChannelMessage t;
        t <- mod_1456.get(0);
        mod_1455.put(1, t);
    endrule
    rule rule_1904;
        ChannelMessage t;
        t <- mod_1469.get(0);
        mod_1470.put(0, t);
    endrule
    rule rule_1905;
        ChannelMessage t;
        t <- mod_1466.get(0);
        mod_1465.put(0, t);
    endrule
    rule rule_1906;
        ChannelMessage t;
        t <- mod_1439.get(0);
        mod_1475.put(0, t);
    endrule
    rule rule_1907;
        ChannelMessage t;
        t <- mod_1447.get(1);
        mod_1448.put(0, t);
    endrule
    rule rule_1908;
        ChannelMessage t;
        t <- mod_1469.get(1);
        mod_1444.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1436.put(0, t);
        end
        if (i == 1) begin
            mod_1452.put(0, t);
        end
        if (i == 2) begin
            mod_1458.put(0, t);
        end
        if (i == 3) begin
            mod_1466.put(0, t);
        end
        if (i == 4) begin
            mod_1472.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_1440.get(0);
        end
        if (i == 0) begin
            t <- mod_1440.get(1);
        end
        if (i == 3) begin
            t <- mod_1440.get(2);
        end
        if (i == 2) begin
            t <- mod_1452.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6070 (Operation_IFC);
    Operation_IFC mod_1477_inner <- mkReshape(2, 64);
    Operation_IFC mod_1477 <- mkDebugOperation(mod_1477_inner, "mod_1477");
    Operation_IFC mod_1478_inner <- mkFlatten(1);
    Operation_IFC mod_1478 <- mkDebugOperation(mod_1478_inner, "mod_1478");
    Operation_IFC mod_1479_inner <- mkFlatten(2);
    Operation_IFC mod_1479 <- mkDebugOperation(mod_1479_inner, "mod_1479");
    Operation_IFC mod_1480_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1480 <- mkDebugOperation(mod_1480_inner, "mod_1480");
    Broadcast_IFC#(4) mod_1481_inner <- mkBroadcast(4);
    Operation_IFC mod_1481 <- mkDebugOperation(mod_1481_inner.op, "mod_1481");
    PMU_IFC mod_1482_bufferize <- mkPMU(2);
    Operation_IFC mod_1482_inner = mod_1482_bufferize.operation;
    Operation_IFC mod_1482 <- mkDebugOperation(mod_1482_inner, "mod_1482");
    Broadcast_IFC#(2) mod_1483_inner <- mkBroadcast(2);
    Operation_IFC mod_1483 <- mkDebugOperation(mod_1483_inner.op, "mod_1483");
    PMU_IFC mod_1484_bufferize <- mkPMU(1);
    Operation_IFC mod_1484_inner = mod_1484_bufferize.operation;
    Operation_IFC mod_1484 <- mkDebugOperation(mod_1484_inner, "mod_1484");
    Operation_IFC mod_1485_inner <- mkBinaryMap(1120, matmul_t_tile);
    Operation_IFC mod_1485 <- mkDebugOperation(mod_1485_inner, "mod_1485");
    Operation_IFC mod_1486_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1486 <- mkDebugOperation(mod_1486_inner, "mod_1486");
    Operation_IFC mod_1487_inner <- mkBinaryMap(1888, mul_tile);
    Operation_IFC mod_1487 <- mkDebugOperation(mod_1487_inner, "mod_1487");
    PMU_IFC mod_1488_bufferize <- mkPMU(1);
    Operation_IFC mod_1488_inner = mod_1488_bufferize.operation;
    Operation_IFC mod_1488 <- mkDebugOperation(mod_1488_inner, "mod_1488");
    Operation_IFC mod_1489_inner <- mkBinaryMap(2491, matmul_t_tile);
    Operation_IFC mod_1489 <- mkDebugOperation(mod_1489_inner, "mod_1489");
    Operation_IFC mod_1490_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1490 <- mkDebugOperation(mod_1490_inner, "mod_1490");
    Operation_IFC mod_1491_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1491 <- mkDebugOperation(mod_1491_inner, "mod_1491");
    Operation_IFC mod_1492_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1492 <- mkDebugOperation(mod_1492_inner, "mod_1492");
    Operation_IFC mod_1493_inner <- mkBinaryMap(2787, mul_tile);
    Operation_IFC mod_1493 <- mkDebugOperation(mod_1493_inner, "mod_1493");
    PMU_IFC mod_1494_bufferize <- mkPMU(1);
    Operation_IFC mod_1494_inner = mod_1494_bufferize.operation;
    Operation_IFC mod_1494 <- mkDebugOperation(mod_1494_inner, "mod_1494");
    PMU_IFC mod_1495_bufferize <- mkPMU(2);
    Operation_IFC mod_1495_inner = mod_1495_bufferize.operation;
    Operation_IFC mod_1495 <- mkDebugOperation(mod_1495_inner, "mod_1495");
    PMU_IFC mod_1496_bufferize <- mkPMU(2);
    Operation_IFC mod_1496_inner = mod_1496_bufferize.operation;
    Operation_IFC mod_1496 <- mkDebugOperation(mod_1496_inner, "mod_1496");
    Operation_IFC mod_1497_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1497 <- mkDebugOperation(mod_1497_inner, "mod_1497");
    Operation_IFC mod_1498_inner <- mkFlatten(1);
    Operation_IFC mod_1498 <- mkDebugOperation(mod_1498_inner, "mod_1498");
    Operation_IFC mod_1499_inner <- mkFlatten(0);
    Operation_IFC mod_1499 <- mkDebugOperation(mod_1499_inner, "mod_1499");
    Operation_IFC mod_1500_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1500 <- mkDebugOperation(mod_1500_inner, "mod_1500");
    Operation_IFC mod_1501_inner <- mkUnaryMap(1760, silu_tile);
    Operation_IFC mod_1501 <- mkDebugOperation(mod_1501_inner, "mod_1501");
    Operation_IFC mod_1502_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1502 <- mkDebugOperation(mod_1502_inner, "mod_1502");
    Operation_IFC mod_1503_inner <- mkBinaryMap(1632, matmul_t_tile);
    Operation_IFC mod_1503 <- mkDebugOperation(mod_1503_inner, "mod_1503");
    PMU_IFC mod_1504_bufferize <- mkPMU(2);
    Operation_IFC mod_1504_inner = mod_1504_bufferize.operation;
    Operation_IFC mod_1504 <- mkDebugOperation(mod_1504_inner, "mod_1504");
    Operation_IFC mod_1505_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1505 <- mkDebugOperation(mod_1505_inner, "mod_1505");
    Operation_IFC mod_1506_inner <- mkFlatten(1);
    Operation_IFC mod_1506 <- mkDebugOperation(mod_1506_inner, "mod_1506");
    Operation_IFC mod_1507_inner <- mkFlatten(0);
    Operation_IFC mod_1507 <- mkDebugOperation(mod_1507_inner, "mod_1507");
    PMU_IFC mod_1508_bufferize <- mkPMU(1);
    Operation_IFC mod_1508_inner = mod_1508_bufferize.operation;
    Operation_IFC mod_1508 <- mkDebugOperation(mod_1508_inner, "mod_1508");
    Operation_IFC mod_1509_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1509 <- mkDebugOperation(mod_1509_inner, "mod_1509");
    PMU_IFC mod_1510_bufferize <- mkPMU(2);
    Operation_IFC mod_1510_inner = mod_1510_bufferize.operation;
    Operation_IFC mod_1510 <- mkDebugOperation(mod_1510_inner, "mod_1510");
    Operation_IFC mod_1511_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1511 <- mkDebugOperation(mod_1511_inner, "mod_1511");
    Operation_IFC mod_1512_inner <- mkFlatten(1);
    Operation_IFC mod_1512 <- mkDebugOperation(mod_1512_inner, "mod_1512");
    Operation_IFC mod_1513_inner <- mkFlatten(0);
    Operation_IFC mod_1513 <- mkDebugOperation(mod_1513_inner, "mod_1513");
    Operation_IFC mod_1514_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1514 <- mkDebugOperation(mod_1514_inner, "mod_1514");
    Operation_IFC mod_1515_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1515 <- mkDebugOperation(mod_1515_inner, "mod_1515");
    PMU_IFC mod_1516_bufferize <- mkPMU(2);
    Operation_IFC mod_1516_inner = mod_1516_bufferize.operation;
    Operation_IFC mod_1516 <- mkDebugOperation(mod_1516_inner, "mod_1516");
    rule rule_1909;
        ChannelMessage t;
        t <- mod_1483.get(1);
        mod_1484.put(0, t);
    endrule
    rule rule_1910;
        ChannelMessage t;
        t <- mod_1505.get(0);
        mod_1504.put(1, t);
    endrule
    rule rule_1911;
        ChannelMessage t;
        t <- mod_1496.get(1);
        mod_1489.put(1, t);
    endrule
    rule rule_1912;
        ChannelMessage t;
        t <- mod_1508.get(1);
        mod_1503.put(0, t);
    endrule
    rule rule_1913;
        ChannelMessage t;
        t <- mod_1510.get(0);
        mod_1511.put(0, t);
    endrule
    rule rule_1914;
        ChannelMessage t;
        t <- mod_1486.get(0);
        mod_1487.put(0, t);
    endrule
    rule rule_1915;
        ChannelMessage t;
        t <- mod_1508.get(0);
        mod_1509.put(0, t);
    endrule
    rule rule_1916;
        ChannelMessage t;
        t <- mod_1482.get(1);
        mod_1483.put(0, t);
    endrule
    rule rule_1917;
        ChannelMessage t;
        t <- mod_1481.get(3);
        mod_1482.put(0, t);
    endrule
    rule rule_1918;
        ChannelMessage t;
        t <- mod_1506.get(0);
        mod_1504.put(0, t);
    endrule
    rule rule_1919;
        ChannelMessage t;
        t <- mod_1514.get(0);
        mod_1484.put(1, t);
    endrule
    rule rule_1920;
        ChannelMessage t;
        t <- mod_1484.get(1);
        mod_1485.put(0, t);
    endrule
    rule rule_1921;
        ChannelMessage t;
        t <- mod_1492.get(0);
        mod_1494.put(0, t);
    endrule
    rule rule_1922;
        ChannelMessage t;
        t <- mod_1492.get(1);
        mod_1493.put(1, t);
    endrule
    rule rule_1923;
        ChannelMessage t;
        t <- mod_1495.get(1);
        mod_1491.put(1, t);
    endrule
    rule rule_1924;
        ChannelMessage t;
        t <- mod_1515.get(0);
        mod_1482.put(1, t);
    endrule
    rule rule_1925;
        ChannelMessage t;
        t <- mod_1509.get(0);
        mod_1508.put(1, t);
    endrule
    rule rule_1926;
        ChannelMessage t;
        t <- mod_1477.get(0);
        mod_1478.put(0, t);
    endrule
    rule rule_1927;
        ChannelMessage t;
        t <- mod_1482.get(0);
        mod_1515.put(0, t);
    endrule
    rule rule_1928;
        ChannelMessage t;
        t <- mod_1507.get(0);
        mod_1506.put(0, t);
    endrule
    rule rule_1929;
        ChannelMessage t;
        t <- mod_1485.get(0);
        mod_1486.put(0, t);
    endrule
    rule rule_1930;
        ChannelMessage t;
        t <- mod_1484.get(0);
        mod_1514.put(0, t);
    endrule
    rule rule_1931;
        ChannelMessage t;
        t <- mod_1487.get(0);
        mod_1488.put(0, t);
    endrule
    rule rule_1932;
        ChannelMessage t;
        t <- mod_1516.get(0);
        mod_1516.put(1, t);
    endrule
    rule rule_1933;
        ChannelMessage t;
        t <- mod_1500.get(0);
        mod_1488.put(1, t);
    endrule
    rule rule_1934;
        ChannelMessage t;
        t <- mod_1489.get(0);
        mod_1490.put(0, t);
    endrule
    rule rule_1935;
        ChannelMessage t;
        t <- mod_1491.get(1);
        mod_1492.put(0, t);
    endrule
    rule rule_1936;
        ChannelMessage t;
        t <- mod_1488.get(1);
        mod_1489.put(0, t);
    endrule
    rule rule_1937;
        ChannelMessage t;
        t <- mod_1494.get(0);
        mod_1494.put(1, t);
    endrule
    rule rule_1938;
        ChannelMessage t;
        t <- mod_1480.get(0);
        mod_1516.put(0, t);
    endrule
    rule rule_1939;
        ChannelMessage t;
        t <- mod_1478.get(0);
        mod_1479.put(0, t);
    endrule
    rule rule_1940;
        ChannelMessage t;
        t <- mod_1497.get(0);
        mod_1496.put(1, t);
    endrule
    rule rule_1941;
        ChannelMessage t;
        t <- mod_1495.get(0);
        mod_1495.put(1, t);
    endrule
    rule rule_1942;
        ChannelMessage t;
        t <- mod_1490.get(0);
        mod_1491.put(0, t);
    endrule
    rule rule_1943;
        ChannelMessage t;
        t <- mod_1491.get(0);
        mod_1495.put(0, t);
    endrule
    rule rule_1944;
        ChannelMessage t;
        t <- mod_1511.get(0);
        mod_1510.put(1, t);
    endrule
    rule rule_1945;
        ChannelMessage t;
        t <- mod_1501.get(0);
        mod_1487.put(1, t);
    endrule
    rule rule_1946;
        ChannelMessage t;
        t <- mod_1488.get(0);
        mod_1500.put(0, t);
    endrule
    rule rule_1947;
        ChannelMessage t;
        t <- mod_1504.get(0);
        mod_1505.put(0, t);
    endrule
    rule rule_1948;
        ChannelMessage t;
        t <- mod_1483.get(0);
        mod_1508.put(0, t);
    endrule
    rule rule_1949;
        ChannelMessage t;
        t <- mod_1496.get(0);
        mod_1497.put(0, t);
    endrule
    rule rule_1950;
        ChannelMessage t;
        t <- mod_1479.get(0);
        mod_1480.put(0, t);
    endrule
    rule rule_1951;
        ChannelMessage t;
        t <- mod_1504.get(1);
        mod_1503.put(1, t);
    endrule
    rule rule_1952;
        ChannelMessage t;
        t <- mod_1502.get(0);
        mod_1501.put(0, t);
    endrule
    rule rule_1953;
        ChannelMessage t;
        t <- mod_1513.get(0);
        mod_1512.put(0, t);
    endrule
    rule rule_1954;
        ChannelMessage t;
        t <- mod_1510.get(1);
        mod_1485.put(1, t);
    endrule
    rule rule_1955;
        ChannelMessage t;
        t <- mod_1503.get(0);
        mod_1502.put(0, t);
    endrule
    rule rule_1956;
        ChannelMessage t;
        t <- mod_1498.get(0);
        mod_1496.put(0, t);
    endrule
    rule rule_1957;
        ChannelMessage t;
        t <- mod_1480.get(1);
        mod_1481.put(0, t);
    endrule
    rule rule_1958;
        ChannelMessage t;
        t <- mod_1512.get(0);
        mod_1510.put(0, t);
    endrule
    rule rule_1959;
        ChannelMessage t;
        t <- mod_1494.get(1);
        mod_1492.put(1, t);
    endrule
    rule rule_1960;
        ChannelMessage t;
        t <- mod_1499.get(0);
        mod_1498.put(0, t);
    endrule
    rule rule_1961;
        ChannelMessage t;
        t <- mod_1516.get(1);
        mod_1480.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1477.put(0, t);
        end
        if (i == 1) begin
            mod_1493.put(0, t);
        end
        if (i == 2) begin
            mod_1499.put(0, t);
        end
        if (i == 3) begin
            mod_1507.put(0, t);
        end
        if (i == 4) begin
            mod_1513.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_1481.get(0);
        end
        if (i == 1) begin
            t <- mod_1481.get(1);
        end
        if (i == 3) begin
            t <- mod_1481.get(2);
        end
        if (i == 2) begin
            t <- mod_1493.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6071 (Operation_IFC);
    Operation_IFC mod_1518_inner <- mkReshape(2, 64);
    Operation_IFC mod_1518 <- mkDebugOperation(mod_1518_inner, "mod_1518");
    Operation_IFC mod_1519_inner <- mkFlatten(1);
    Operation_IFC mod_1519 <- mkDebugOperation(mod_1519_inner, "mod_1519");
    Operation_IFC mod_1520_inner <- mkFlatten(2);
    Operation_IFC mod_1520 <- mkDebugOperation(mod_1520_inner, "mod_1520");
    Operation_IFC mod_1521_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1521 <- mkDebugOperation(mod_1521_inner, "mod_1521");
    Broadcast_IFC#(4) mod_1522_inner <- mkBroadcast(4);
    Operation_IFC mod_1522 <- mkDebugOperation(mod_1522_inner.op, "mod_1522");
    PMU_IFC mod_1523_bufferize <- mkPMU(2);
    Operation_IFC mod_1523_inner = mod_1523_bufferize.operation;
    Operation_IFC mod_1523 <- mkDebugOperation(mod_1523_inner, "mod_1523");
    Broadcast_IFC#(2) mod_1524_inner <- mkBroadcast(2);
    Operation_IFC mod_1524 <- mkDebugOperation(mod_1524_inner.op, "mod_1524");
    PMU_IFC mod_1525_bufferize <- mkPMU(1);
    Operation_IFC mod_1525_inner = mod_1525_bufferize.operation;
    Operation_IFC mod_1525 <- mkDebugOperation(mod_1525_inner, "mod_1525");
    Operation_IFC mod_1526_inner <- mkBinaryMap(1119, matmul_t_tile);
    Operation_IFC mod_1526 <- mkDebugOperation(mod_1526_inner, "mod_1526");
    Operation_IFC mod_1527_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1527 <- mkDebugOperation(mod_1527_inner, "mod_1527");
    Operation_IFC mod_1528_inner <- mkBinaryMap(1887, mul_tile);
    Operation_IFC mod_1528 <- mkDebugOperation(mod_1528_inner, "mod_1528");
    PMU_IFC mod_1529_bufferize <- mkPMU(1);
    Operation_IFC mod_1529_inner = mod_1529_bufferize.operation;
    Operation_IFC mod_1529 <- mkDebugOperation(mod_1529_inner, "mod_1529");
    Operation_IFC mod_1530_inner <- mkBinaryMap(2489, matmul_t_tile);
    Operation_IFC mod_1530 <- mkDebugOperation(mod_1530_inner, "mod_1530");
    Operation_IFC mod_1531_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1531 <- mkDebugOperation(mod_1531_inner, "mod_1531");
    Operation_IFC mod_1532_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1532 <- mkDebugOperation(mod_1532_inner, "mod_1532");
    Operation_IFC mod_1533_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1533 <- mkDebugOperation(mod_1533_inner, "mod_1533");
    Operation_IFC mod_1534_inner <- mkBinaryMap(2786, mul_tile);
    Operation_IFC mod_1534 <- mkDebugOperation(mod_1534_inner, "mod_1534");
    PMU_IFC mod_1535_bufferize <- mkPMU(1);
    Operation_IFC mod_1535_inner = mod_1535_bufferize.operation;
    Operation_IFC mod_1535 <- mkDebugOperation(mod_1535_inner, "mod_1535");
    PMU_IFC mod_1536_bufferize <- mkPMU(2);
    Operation_IFC mod_1536_inner = mod_1536_bufferize.operation;
    Operation_IFC mod_1536 <- mkDebugOperation(mod_1536_inner, "mod_1536");
    PMU_IFC mod_1537_bufferize <- mkPMU(2);
    Operation_IFC mod_1537_inner = mod_1537_bufferize.operation;
    Operation_IFC mod_1537 <- mkDebugOperation(mod_1537_inner, "mod_1537");
    Operation_IFC mod_1538_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1538 <- mkDebugOperation(mod_1538_inner, "mod_1538");
    Operation_IFC mod_1539_inner <- mkFlatten(1);
    Operation_IFC mod_1539 <- mkDebugOperation(mod_1539_inner, "mod_1539");
    Operation_IFC mod_1540_inner <- mkFlatten(0);
    Operation_IFC mod_1540 <- mkDebugOperation(mod_1540_inner, "mod_1540");
    Operation_IFC mod_1541_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1541 <- mkDebugOperation(mod_1541_inner, "mod_1541");
    Operation_IFC mod_1542_inner <- mkUnaryMap(1759, silu_tile);
    Operation_IFC mod_1542 <- mkDebugOperation(mod_1542_inner, "mod_1542");
    Operation_IFC mod_1543_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1543 <- mkDebugOperation(mod_1543_inner, "mod_1543");
    Operation_IFC mod_1544_inner <- mkBinaryMap(1631, matmul_t_tile);
    Operation_IFC mod_1544 <- mkDebugOperation(mod_1544_inner, "mod_1544");
    PMU_IFC mod_1545_bufferize <- mkPMU(2);
    Operation_IFC mod_1545_inner = mod_1545_bufferize.operation;
    Operation_IFC mod_1545 <- mkDebugOperation(mod_1545_inner, "mod_1545");
    Operation_IFC mod_1546_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1546 <- mkDebugOperation(mod_1546_inner, "mod_1546");
    Operation_IFC mod_1547_inner <- mkFlatten(1);
    Operation_IFC mod_1547 <- mkDebugOperation(mod_1547_inner, "mod_1547");
    Operation_IFC mod_1548_inner <- mkFlatten(0);
    Operation_IFC mod_1548 <- mkDebugOperation(mod_1548_inner, "mod_1548");
    PMU_IFC mod_1549_bufferize <- mkPMU(1);
    Operation_IFC mod_1549_inner = mod_1549_bufferize.operation;
    Operation_IFC mod_1549 <- mkDebugOperation(mod_1549_inner, "mod_1549");
    Operation_IFC mod_1550_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1550 <- mkDebugOperation(mod_1550_inner, "mod_1550");
    PMU_IFC mod_1551_bufferize <- mkPMU(2);
    Operation_IFC mod_1551_inner = mod_1551_bufferize.operation;
    Operation_IFC mod_1551 <- mkDebugOperation(mod_1551_inner, "mod_1551");
    Operation_IFC mod_1552_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1552 <- mkDebugOperation(mod_1552_inner, "mod_1552");
    Operation_IFC mod_1553_inner <- mkFlatten(1);
    Operation_IFC mod_1553 <- mkDebugOperation(mod_1553_inner, "mod_1553");
    Operation_IFC mod_1554_inner <- mkFlatten(0);
    Operation_IFC mod_1554 <- mkDebugOperation(mod_1554_inner, "mod_1554");
    Operation_IFC mod_1555_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1555 <- mkDebugOperation(mod_1555_inner, "mod_1555");
    Operation_IFC mod_1556_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1556 <- mkDebugOperation(mod_1556_inner, "mod_1556");
    PMU_IFC mod_1557_bufferize <- mkPMU(2);
    Operation_IFC mod_1557_inner = mod_1557_bufferize.operation;
    Operation_IFC mod_1557 <- mkDebugOperation(mod_1557_inner, "mod_1557");
    rule rule_1962;
        ChannelMessage t;
        t <- mod_1549.get(0);
        mod_1550.put(0, t);
    endrule
    rule rule_1963;
        ChannelMessage t;
        t <- mod_1525.get(1);
        mod_1526.put(0, t);
    endrule
    rule rule_1964;
        ChannelMessage t;
        t <- mod_1550.get(0);
        mod_1549.put(1, t);
    endrule
    rule rule_1965;
        ChannelMessage t;
        t <- mod_1551.get(1);
        mod_1526.put(1, t);
    endrule
    rule rule_1966;
        ChannelMessage t;
        t <- mod_1552.get(0);
        mod_1551.put(1, t);
    endrule
    rule rule_1967;
        ChannelMessage t;
        t <- mod_1553.get(0);
        mod_1551.put(0, t);
    endrule
    rule rule_1968;
        ChannelMessage t;
        t <- mod_1535.get(1);
        mod_1533.put(1, t);
    endrule
    rule rule_1969;
        ChannelMessage t;
        t <- mod_1521.get(1);
        mod_1522.put(0, t);
    endrule
    rule rule_1970;
        ChannelMessage t;
        t <- mod_1545.get(0);
        mod_1546.put(0, t);
    endrule
    rule rule_1971;
        ChannelMessage t;
        t <- mod_1548.get(0);
        mod_1547.put(0, t);
    endrule
    rule rule_1972;
        ChannelMessage t;
        t <- mod_1529.get(1);
        mod_1530.put(0, t);
    endrule
    rule rule_1973;
        ChannelMessage t;
        t <- mod_1524.get(0);
        mod_1549.put(0, t);
    endrule
    rule rule_1974;
        ChannelMessage t;
        t <- mod_1555.get(0);
        mod_1525.put(1, t);
    endrule
    rule rule_1975;
        ChannelMessage t;
        t <- mod_1521.get(0);
        mod_1557.put(0, t);
    endrule
    rule rule_1976;
        ChannelMessage t;
        t <- mod_1528.get(0);
        mod_1529.put(0, t);
    endrule
    rule rule_1977;
        ChannelMessage t;
        t <- mod_1556.get(0);
        mod_1523.put(1, t);
    endrule
    rule rule_1978;
        ChannelMessage t;
        t <- mod_1549.get(1);
        mod_1544.put(0, t);
    endrule
    rule rule_1979;
        ChannelMessage t;
        t <- mod_1530.get(0);
        mod_1531.put(0, t);
    endrule
    rule rule_1980;
        ChannelMessage t;
        t <- mod_1543.get(0);
        mod_1542.put(0, t);
    endrule
    rule rule_1981;
        ChannelMessage t;
        t <- mod_1532.get(1);
        mod_1533.put(0, t);
    endrule
    rule rule_1982;
        ChannelMessage t;
        t <- mod_1542.get(0);
        mod_1528.put(1, t);
    endrule
    rule rule_1983;
        ChannelMessage t;
        t <- mod_1537.get(1);
        mod_1530.put(1, t);
    endrule
    rule rule_1984;
        ChannelMessage t;
        t <- mod_1529.get(0);
        mod_1541.put(0, t);
    endrule
    rule rule_1985;
        ChannelMessage t;
        t <- mod_1526.get(0);
        mod_1527.put(0, t);
    endrule
    rule rule_1986;
        ChannelMessage t;
        t <- mod_1531.get(0);
        mod_1532.put(0, t);
    endrule
    rule rule_1987;
        ChannelMessage t;
        t <- mod_1533.get(0);
        mod_1535.put(0, t);
    endrule
    rule rule_1988;
        ChannelMessage t;
        t <- mod_1537.get(0);
        mod_1538.put(0, t);
    endrule
    rule rule_1989;
        ChannelMessage t;
        t <- mod_1540.get(0);
        mod_1539.put(0, t);
    endrule
    rule rule_1990;
        ChannelMessage t;
        t <- mod_1536.get(1);
        mod_1532.put(1, t);
    endrule
    rule rule_1991;
        ChannelMessage t;
        t <- mod_1545.get(1);
        mod_1544.put(1, t);
    endrule
    rule rule_1992;
        ChannelMessage t;
        t <- mod_1535.get(0);
        mod_1535.put(1, t);
    endrule
    rule rule_1993;
        ChannelMessage t;
        t <- mod_1539.get(0);
        mod_1537.put(0, t);
    endrule
    rule rule_1994;
        ChannelMessage t;
        t <- mod_1546.get(0);
        mod_1545.put(1, t);
    endrule
    rule rule_1995;
        ChannelMessage t;
        t <- mod_1557.get(0);
        mod_1557.put(1, t);
    endrule
    rule rule_1996;
        ChannelMessage t;
        t <- mod_1541.get(0);
        mod_1529.put(1, t);
    endrule
    rule rule_1997;
        ChannelMessage t;
        t <- mod_1527.get(0);
        mod_1528.put(0, t);
    endrule
    rule rule_1998;
        ChannelMessage t;
        t <- mod_1519.get(0);
        mod_1520.put(0, t);
    endrule
    rule rule_1999;
        ChannelMessage t;
        t <- mod_1525.get(0);
        mod_1555.put(0, t);
    endrule
    rule rule_2000;
        ChannelMessage t;
        t <- mod_1547.get(0);
        mod_1545.put(0, t);
    endrule
    rule rule_2001;
        ChannelMessage t;
        t <- mod_1522.get(3);
        mod_1523.put(0, t);
    endrule
    rule rule_2002;
        ChannelMessage t;
        t <- mod_1524.get(1);
        mod_1525.put(0, t);
    endrule
    rule rule_2003;
        ChannelMessage t;
        t <- mod_1523.get(1);
        mod_1524.put(0, t);
    endrule
    rule rule_2004;
        ChannelMessage t;
        t <- mod_1523.get(0);
        mod_1556.put(0, t);
    endrule
    rule rule_2005;
        ChannelMessage t;
        t <- mod_1532.get(0);
        mod_1536.put(0, t);
    endrule
    rule rule_2006;
        ChannelMessage t;
        t <- mod_1544.get(0);
        mod_1543.put(0, t);
    endrule
    rule rule_2007;
        ChannelMessage t;
        t <- mod_1533.get(1);
        mod_1534.put(1, t);
    endrule
    rule rule_2008;
        ChannelMessage t;
        t <- mod_1536.get(0);
        mod_1536.put(1, t);
    endrule
    rule rule_2009;
        ChannelMessage t;
        t <- mod_1551.get(0);
        mod_1552.put(0, t);
    endrule
    rule rule_2010;
        ChannelMessage t;
        t <- mod_1557.get(1);
        mod_1521.put(1, t);
    endrule
    rule rule_2011;
        ChannelMessage t;
        t <- mod_1518.get(0);
        mod_1519.put(0, t);
    endrule
    rule rule_2012;
        ChannelMessage t;
        t <- mod_1554.get(0);
        mod_1553.put(0, t);
    endrule
    rule rule_2013;
        ChannelMessage t;
        t <- mod_1520.get(0);
        mod_1521.put(0, t);
    endrule
    rule rule_2014;
        ChannelMessage t;
        t <- mod_1538.get(0);
        mod_1537.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1518.put(0, t);
        end
        if (i == 1) begin
            mod_1534.put(0, t);
        end
        if (i == 2) begin
            mod_1540.put(0, t);
        end
        if (i == 3) begin
            mod_1548.put(0, t);
        end
        if (i == 4) begin
            mod_1554.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 2) begin
            t <- mod_1522.get(0);
        end
        if (i == 0) begin
            t <- mod_1522.get(1);
        end
        if (i == 3) begin
            t <- mod_1522.get(2);
        end
        if (i == 1) begin
            t <- mod_1534.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6072 (Operation_IFC);
    Operation_IFC mod_1559_inner <- mkReshape(2, 64);
    Operation_IFC mod_1559 <- mkDebugOperation(mod_1559_inner, "mod_1559");
    Operation_IFC mod_1560_inner <- mkFlatten(1);
    Operation_IFC mod_1560 <- mkDebugOperation(mod_1560_inner, "mod_1560");
    Operation_IFC mod_1561_inner <- mkFlatten(2);
    Operation_IFC mod_1561 <- mkDebugOperation(mod_1561_inner, "mod_1561");
    Operation_IFC mod_1562_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1562 <- mkDebugOperation(mod_1562_inner, "mod_1562");
    Broadcast_IFC#(4) mod_1563_inner <- mkBroadcast(4);
    Operation_IFC mod_1563 <- mkDebugOperation(mod_1563_inner.op, "mod_1563");
    PMU_IFC mod_1564_bufferize <- mkPMU(2);
    Operation_IFC mod_1564_inner = mod_1564_bufferize.operation;
    Operation_IFC mod_1564 <- mkDebugOperation(mod_1564_inner, "mod_1564");
    Broadcast_IFC#(2) mod_1565_inner <- mkBroadcast(2);
    Operation_IFC mod_1565 <- mkDebugOperation(mod_1565_inner.op, "mod_1565");
    PMU_IFC mod_1566_bufferize <- mkPMU(1);
    Operation_IFC mod_1566_inner = mod_1566_bufferize.operation;
    Operation_IFC mod_1566 <- mkDebugOperation(mod_1566_inner, "mod_1566");
    Operation_IFC mod_1567_inner <- mkBinaryMap(1118, matmul_t_tile);
    Operation_IFC mod_1567 <- mkDebugOperation(mod_1567_inner, "mod_1567");
    Operation_IFC mod_1568_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1568 <- mkDebugOperation(mod_1568_inner, "mod_1568");
    Operation_IFC mod_1569_inner <- mkBinaryMap(1886, mul_tile);
    Operation_IFC mod_1569 <- mkDebugOperation(mod_1569_inner, "mod_1569");
    PMU_IFC mod_1570_bufferize <- mkPMU(1);
    Operation_IFC mod_1570_inner = mod_1570_bufferize.operation;
    Operation_IFC mod_1570 <- mkDebugOperation(mod_1570_inner, "mod_1570");
    Operation_IFC mod_1571_inner <- mkBinaryMap(2487, matmul_t_tile);
    Operation_IFC mod_1571 <- mkDebugOperation(mod_1571_inner, "mod_1571");
    Operation_IFC mod_1572_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1572 <- mkDebugOperation(mod_1572_inner, "mod_1572");
    Operation_IFC mod_1573_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1573 <- mkDebugOperation(mod_1573_inner, "mod_1573");
    Operation_IFC mod_1574_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1574 <- mkDebugOperation(mod_1574_inner, "mod_1574");
    Operation_IFC mod_1575_inner <- mkBinaryMap(2785, mul_tile);
    Operation_IFC mod_1575 <- mkDebugOperation(mod_1575_inner, "mod_1575");
    PMU_IFC mod_1576_bufferize <- mkPMU(1);
    Operation_IFC mod_1576_inner = mod_1576_bufferize.operation;
    Operation_IFC mod_1576 <- mkDebugOperation(mod_1576_inner, "mod_1576");
    PMU_IFC mod_1577_bufferize <- mkPMU(2);
    Operation_IFC mod_1577_inner = mod_1577_bufferize.operation;
    Operation_IFC mod_1577 <- mkDebugOperation(mod_1577_inner, "mod_1577");
    PMU_IFC mod_1578_bufferize <- mkPMU(2);
    Operation_IFC mod_1578_inner = mod_1578_bufferize.operation;
    Operation_IFC mod_1578 <- mkDebugOperation(mod_1578_inner, "mod_1578");
    Operation_IFC mod_1579_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1579 <- mkDebugOperation(mod_1579_inner, "mod_1579");
    Operation_IFC mod_1580_inner <- mkFlatten(1);
    Operation_IFC mod_1580 <- mkDebugOperation(mod_1580_inner, "mod_1580");
    Operation_IFC mod_1581_inner <- mkFlatten(0);
    Operation_IFC mod_1581 <- mkDebugOperation(mod_1581_inner, "mod_1581");
    Operation_IFC mod_1582_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1582 <- mkDebugOperation(mod_1582_inner, "mod_1582");
    Operation_IFC mod_1583_inner <- mkUnaryMap(1758, silu_tile);
    Operation_IFC mod_1583 <- mkDebugOperation(mod_1583_inner, "mod_1583");
    Operation_IFC mod_1584_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1584 <- mkDebugOperation(mod_1584_inner, "mod_1584");
    Operation_IFC mod_1585_inner <- mkBinaryMap(1630, matmul_t_tile);
    Operation_IFC mod_1585 <- mkDebugOperation(mod_1585_inner, "mod_1585");
    PMU_IFC mod_1586_bufferize <- mkPMU(2);
    Operation_IFC mod_1586_inner = mod_1586_bufferize.operation;
    Operation_IFC mod_1586 <- mkDebugOperation(mod_1586_inner, "mod_1586");
    Operation_IFC mod_1587_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1587 <- mkDebugOperation(mod_1587_inner, "mod_1587");
    Operation_IFC mod_1588_inner <- mkFlatten(1);
    Operation_IFC mod_1588 <- mkDebugOperation(mod_1588_inner, "mod_1588");
    Operation_IFC mod_1589_inner <- mkFlatten(0);
    Operation_IFC mod_1589 <- mkDebugOperation(mod_1589_inner, "mod_1589");
    PMU_IFC mod_1590_bufferize <- mkPMU(1);
    Operation_IFC mod_1590_inner = mod_1590_bufferize.operation;
    Operation_IFC mod_1590 <- mkDebugOperation(mod_1590_inner, "mod_1590");
    Operation_IFC mod_1591_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1591 <- mkDebugOperation(mod_1591_inner, "mod_1591");
    PMU_IFC mod_1592_bufferize <- mkPMU(2);
    Operation_IFC mod_1592_inner = mod_1592_bufferize.operation;
    Operation_IFC mod_1592 <- mkDebugOperation(mod_1592_inner, "mod_1592");
    Operation_IFC mod_1593_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1593 <- mkDebugOperation(mod_1593_inner, "mod_1593");
    Operation_IFC mod_1594_inner <- mkFlatten(1);
    Operation_IFC mod_1594 <- mkDebugOperation(mod_1594_inner, "mod_1594");
    Operation_IFC mod_1595_inner <- mkFlatten(0);
    Operation_IFC mod_1595 <- mkDebugOperation(mod_1595_inner, "mod_1595");
    Operation_IFC mod_1596_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1596 <- mkDebugOperation(mod_1596_inner, "mod_1596");
    Operation_IFC mod_1597_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1597 <- mkDebugOperation(mod_1597_inner, "mod_1597");
    PMU_IFC mod_1598_bufferize <- mkPMU(2);
    Operation_IFC mod_1598_inner = mod_1598_bufferize.operation;
    Operation_IFC mod_1598 <- mkDebugOperation(mod_1598_inner, "mod_1598");
    rule rule_2015;
        ChannelMessage t;
        t <- mod_1590.get(0);
        mod_1591.put(0, t);
    endrule
    rule rule_2016;
        ChannelMessage t;
        t <- mod_1597.get(0);
        mod_1564.put(1, t);
    endrule
    rule rule_2017;
        ChannelMessage t;
        t <- mod_1577.get(1);
        mod_1573.put(1, t);
    endrule
    rule rule_2018;
        ChannelMessage t;
        t <- mod_1585.get(0);
        mod_1584.put(0, t);
    endrule
    rule rule_2019;
        ChannelMessage t;
        t <- mod_1566.get(0);
        mod_1596.put(0, t);
    endrule
    rule rule_2020;
        ChannelMessage t;
        t <- mod_1561.get(0);
        mod_1562.put(0, t);
    endrule
    rule rule_2021;
        ChannelMessage t;
        t <- mod_1559.get(0);
        mod_1560.put(0, t);
    endrule
    rule rule_2022;
        ChannelMessage t;
        t <- mod_1564.get(1);
        mod_1565.put(0, t);
    endrule
    rule rule_2023;
        ChannelMessage t;
        t <- mod_1567.get(0);
        mod_1568.put(0, t);
    endrule
    rule rule_2024;
        ChannelMessage t;
        t <- mod_1577.get(0);
        mod_1577.put(1, t);
    endrule
    rule rule_2025;
        ChannelMessage t;
        t <- mod_1592.get(1);
        mod_1567.put(1, t);
    endrule
    rule rule_2026;
        ChannelMessage t;
        t <- mod_1581.get(0);
        mod_1580.put(0, t);
    endrule
    rule rule_2027;
        ChannelMessage t;
        t <- mod_1586.get(0);
        mod_1587.put(0, t);
    endrule
    rule rule_2028;
        ChannelMessage t;
        t <- mod_1574.get(0);
        mod_1576.put(0, t);
    endrule
    rule rule_2029;
        ChannelMessage t;
        t <- mod_1580.get(0);
        mod_1578.put(0, t);
    endrule
    rule rule_2030;
        ChannelMessage t;
        t <- mod_1562.get(1);
        mod_1563.put(0, t);
    endrule
    rule rule_2031;
        ChannelMessage t;
        t <- mod_1582.get(0);
        mod_1570.put(1, t);
    endrule
    rule rule_2032;
        ChannelMessage t;
        t <- mod_1592.get(0);
        mod_1593.put(0, t);
    endrule
    rule rule_2033;
        ChannelMessage t;
        t <- mod_1598.get(1);
        mod_1562.put(1, t);
    endrule
    rule rule_2034;
        ChannelMessage t;
        t <- mod_1586.get(1);
        mod_1585.put(1, t);
    endrule
    rule rule_2035;
        ChannelMessage t;
        t <- mod_1589.get(0);
        mod_1588.put(0, t);
    endrule
    rule rule_2036;
        ChannelMessage t;
        t <- mod_1560.get(0);
        mod_1561.put(0, t);
    endrule
    rule rule_2037;
        ChannelMessage t;
        t <- mod_1591.get(0);
        mod_1590.put(1, t);
    endrule
    rule rule_2038;
        ChannelMessage t;
        t <- mod_1573.get(0);
        mod_1577.put(0, t);
    endrule
    rule rule_2039;
        ChannelMessage t;
        t <- mod_1590.get(1);
        mod_1585.put(0, t);
    endrule
    rule rule_2040;
        ChannelMessage t;
        t <- mod_1576.get(0);
        mod_1576.put(1, t);
    endrule
    rule rule_2041;
        ChannelMessage t;
        t <- mod_1565.get(1);
        mod_1566.put(0, t);
    endrule
    rule rule_2042;
        ChannelMessage t;
        t <- mod_1573.get(1);
        mod_1574.put(0, t);
    endrule
    rule rule_2043;
        ChannelMessage t;
        t <- mod_1576.get(1);
        mod_1574.put(1, t);
    endrule
    rule rule_2044;
        ChannelMessage t;
        t <- mod_1564.get(0);
        mod_1597.put(0, t);
    endrule
    rule rule_2045;
        ChannelMessage t;
        t <- mod_1578.get(0);
        mod_1579.put(0, t);
    endrule
    rule rule_2046;
        ChannelMessage t;
        t <- mod_1593.get(0);
        mod_1592.put(1, t);
    endrule
    rule rule_2047;
        ChannelMessage t;
        t <- mod_1588.get(0);
        mod_1586.put(0, t);
    endrule
    rule rule_2048;
        ChannelMessage t;
        t <- mod_1566.get(1);
        mod_1567.put(0, t);
    endrule
    rule rule_2049;
        ChannelMessage t;
        t <- mod_1569.get(0);
        mod_1570.put(0, t);
    endrule
    rule rule_2050;
        ChannelMessage t;
        t <- mod_1570.get(1);
        mod_1571.put(0, t);
    endrule
    rule rule_2051;
        ChannelMessage t;
        t <- mod_1596.get(0);
        mod_1566.put(1, t);
    endrule
    rule rule_2052;
        ChannelMessage t;
        t <- mod_1565.get(0);
        mod_1590.put(0, t);
    endrule
    rule rule_2053;
        ChannelMessage t;
        t <- mod_1578.get(1);
        mod_1571.put(1, t);
    endrule
    rule rule_2054;
        ChannelMessage t;
        t <- mod_1584.get(0);
        mod_1583.put(0, t);
    endrule
    rule rule_2055;
        ChannelMessage t;
        t <- mod_1563.get(3);
        mod_1564.put(0, t);
    endrule
    rule rule_2056;
        ChannelMessage t;
        t <- mod_1572.get(0);
        mod_1573.put(0, t);
    endrule
    rule rule_2057;
        ChannelMessage t;
        t <- mod_1570.get(0);
        mod_1582.put(0, t);
    endrule
    rule rule_2058;
        ChannelMessage t;
        t <- mod_1562.get(0);
        mod_1598.put(0, t);
    endrule
    rule rule_2059;
        ChannelMessage t;
        t <- mod_1587.get(0);
        mod_1586.put(1, t);
    endrule
    rule rule_2060;
        ChannelMessage t;
        t <- mod_1594.get(0);
        mod_1592.put(0, t);
    endrule
    rule rule_2061;
        ChannelMessage t;
        t <- mod_1574.get(1);
        mod_1575.put(1, t);
    endrule
    rule rule_2062;
        ChannelMessage t;
        t <- mod_1583.get(0);
        mod_1569.put(1, t);
    endrule
    rule rule_2063;
        ChannelMessage t;
        t <- mod_1568.get(0);
        mod_1569.put(0, t);
    endrule
    rule rule_2064;
        ChannelMessage t;
        t <- mod_1579.get(0);
        mod_1578.put(1, t);
    endrule
    rule rule_2065;
        ChannelMessage t;
        t <- mod_1571.get(0);
        mod_1572.put(0, t);
    endrule
    rule rule_2066;
        ChannelMessage t;
        t <- mod_1595.get(0);
        mod_1594.put(0, t);
    endrule
    rule rule_2067;
        ChannelMessage t;
        t <- mod_1598.get(0);
        mod_1598.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1559.put(0, t);
        end
        if (i == 1) begin
            mod_1575.put(0, t);
        end
        if (i == 2) begin
            mod_1581.put(0, t);
        end
        if (i == 3) begin
            mod_1589.put(0, t);
        end
        if (i == 4) begin
            mod_1595.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_1563.get(0);
        end
        if (i == 0) begin
            t <- mod_1563.get(1);
        end
        if (i == 2) begin
            t <- mod_1563.get(2);
        end
        if (i == 1) begin
            t <- mod_1575.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6073 (Operation_IFC);
    Operation_IFC mod_1600_inner <- mkReshape(2, 64);
    Operation_IFC mod_1600 <- mkDebugOperation(mod_1600_inner, "mod_1600");
    Operation_IFC mod_1601_inner <- mkFlatten(1);
    Operation_IFC mod_1601 <- mkDebugOperation(mod_1601_inner, "mod_1601");
    Operation_IFC mod_1602_inner <- mkFlatten(2);
    Operation_IFC mod_1602 <- mkDebugOperation(mod_1602_inner, "mod_1602");
    Operation_IFC mod_1603_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1603 <- mkDebugOperation(mod_1603_inner, "mod_1603");
    Broadcast_IFC#(4) mod_1604_inner <- mkBroadcast(4);
    Operation_IFC mod_1604 <- mkDebugOperation(mod_1604_inner.op, "mod_1604");
    PMU_IFC mod_1605_bufferize <- mkPMU(2);
    Operation_IFC mod_1605_inner = mod_1605_bufferize.operation;
    Operation_IFC mod_1605 <- mkDebugOperation(mod_1605_inner, "mod_1605");
    Broadcast_IFC#(2) mod_1606_inner <- mkBroadcast(2);
    Operation_IFC mod_1606 <- mkDebugOperation(mod_1606_inner.op, "mod_1606");
    PMU_IFC mod_1607_bufferize <- mkPMU(1);
    Operation_IFC mod_1607_inner = mod_1607_bufferize.operation;
    Operation_IFC mod_1607 <- mkDebugOperation(mod_1607_inner, "mod_1607");
    Operation_IFC mod_1608_inner <- mkBinaryMap(1117, matmul_t_tile);
    Operation_IFC mod_1608 <- mkDebugOperation(mod_1608_inner, "mod_1608");
    Operation_IFC mod_1609_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1609 <- mkDebugOperation(mod_1609_inner, "mod_1609");
    Operation_IFC mod_1610_inner <- mkBinaryMap(1885, mul_tile);
    Operation_IFC mod_1610 <- mkDebugOperation(mod_1610_inner, "mod_1610");
    PMU_IFC mod_1611_bufferize <- mkPMU(1);
    Operation_IFC mod_1611_inner = mod_1611_bufferize.operation;
    Operation_IFC mod_1611 <- mkDebugOperation(mod_1611_inner, "mod_1611");
    Operation_IFC mod_1612_inner <- mkBinaryMap(2485, matmul_t_tile);
    Operation_IFC mod_1612 <- mkDebugOperation(mod_1612_inner, "mod_1612");
    Operation_IFC mod_1613_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1613 <- mkDebugOperation(mod_1613_inner, "mod_1613");
    Operation_IFC mod_1614_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1614 <- mkDebugOperation(mod_1614_inner, "mod_1614");
    Operation_IFC mod_1615_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1615 <- mkDebugOperation(mod_1615_inner, "mod_1615");
    Operation_IFC mod_1616_inner <- mkBinaryMap(2784, mul_tile);
    Operation_IFC mod_1616 <- mkDebugOperation(mod_1616_inner, "mod_1616");
    PMU_IFC mod_1617_bufferize <- mkPMU(1);
    Operation_IFC mod_1617_inner = mod_1617_bufferize.operation;
    Operation_IFC mod_1617 <- mkDebugOperation(mod_1617_inner, "mod_1617");
    PMU_IFC mod_1618_bufferize <- mkPMU(2);
    Operation_IFC mod_1618_inner = mod_1618_bufferize.operation;
    Operation_IFC mod_1618 <- mkDebugOperation(mod_1618_inner, "mod_1618");
    PMU_IFC mod_1619_bufferize <- mkPMU(2);
    Operation_IFC mod_1619_inner = mod_1619_bufferize.operation;
    Operation_IFC mod_1619 <- mkDebugOperation(mod_1619_inner, "mod_1619");
    Operation_IFC mod_1620_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1620 <- mkDebugOperation(mod_1620_inner, "mod_1620");
    Operation_IFC mod_1621_inner <- mkFlatten(1);
    Operation_IFC mod_1621 <- mkDebugOperation(mod_1621_inner, "mod_1621");
    Operation_IFC mod_1622_inner <- mkFlatten(0);
    Operation_IFC mod_1622 <- mkDebugOperation(mod_1622_inner, "mod_1622");
    Operation_IFC mod_1623_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1623 <- mkDebugOperation(mod_1623_inner, "mod_1623");
    Operation_IFC mod_1624_inner <- mkUnaryMap(1757, silu_tile);
    Operation_IFC mod_1624 <- mkDebugOperation(mod_1624_inner, "mod_1624");
    Operation_IFC mod_1625_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1625 <- mkDebugOperation(mod_1625_inner, "mod_1625");
    Operation_IFC mod_1626_inner <- mkBinaryMap(1629, matmul_t_tile);
    Operation_IFC mod_1626 <- mkDebugOperation(mod_1626_inner, "mod_1626");
    PMU_IFC mod_1627_bufferize <- mkPMU(2);
    Operation_IFC mod_1627_inner = mod_1627_bufferize.operation;
    Operation_IFC mod_1627 <- mkDebugOperation(mod_1627_inner, "mod_1627");
    Operation_IFC mod_1628_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1628 <- mkDebugOperation(mod_1628_inner, "mod_1628");
    Operation_IFC mod_1629_inner <- mkFlatten(1);
    Operation_IFC mod_1629 <- mkDebugOperation(mod_1629_inner, "mod_1629");
    Operation_IFC mod_1630_inner <- mkFlatten(0);
    Operation_IFC mod_1630 <- mkDebugOperation(mod_1630_inner, "mod_1630");
    PMU_IFC mod_1631_bufferize <- mkPMU(1);
    Operation_IFC mod_1631_inner = mod_1631_bufferize.operation;
    Operation_IFC mod_1631 <- mkDebugOperation(mod_1631_inner, "mod_1631");
    Operation_IFC mod_1632_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1632 <- mkDebugOperation(mod_1632_inner, "mod_1632");
    PMU_IFC mod_1633_bufferize <- mkPMU(2);
    Operation_IFC mod_1633_inner = mod_1633_bufferize.operation;
    Operation_IFC mod_1633 <- mkDebugOperation(mod_1633_inner, "mod_1633");
    Operation_IFC mod_1634_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1634 <- mkDebugOperation(mod_1634_inner, "mod_1634");
    Operation_IFC mod_1635_inner <- mkFlatten(1);
    Operation_IFC mod_1635 <- mkDebugOperation(mod_1635_inner, "mod_1635");
    Operation_IFC mod_1636_inner <- mkFlatten(0);
    Operation_IFC mod_1636 <- mkDebugOperation(mod_1636_inner, "mod_1636");
    Operation_IFC mod_1637_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1637 <- mkDebugOperation(mod_1637_inner, "mod_1637");
    Operation_IFC mod_1638_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1638 <- mkDebugOperation(mod_1638_inner, "mod_1638");
    PMU_IFC mod_1639_bufferize <- mkPMU(2);
    Operation_IFC mod_1639_inner = mod_1639_bufferize.operation;
    Operation_IFC mod_1639 <- mkDebugOperation(mod_1639_inner, "mod_1639");
    rule rule_2068;
        ChannelMessage t;
        t <- mod_1619.get(0);
        mod_1620.put(0, t);
    endrule
    rule rule_2069;
        ChannelMessage t;
        t <- mod_1613.get(0);
        mod_1614.put(0, t);
    endrule
    rule rule_2070;
        ChannelMessage t;
        t <- mod_1615.get(0);
        mod_1617.put(0, t);
    endrule
    rule rule_2071;
        ChannelMessage t;
        t <- mod_1614.get(0);
        mod_1618.put(0, t);
    endrule
    rule rule_2072;
        ChannelMessage t;
        t <- mod_1611.get(0);
        mod_1623.put(0, t);
    endrule
    rule rule_2073;
        ChannelMessage t;
        t <- mod_1618.get(1);
        mod_1614.put(1, t);
    endrule
    rule rule_2074;
        ChannelMessage t;
        t <- mod_1612.get(0);
        mod_1613.put(0, t);
    endrule
    rule rule_2075;
        ChannelMessage t;
        t <- mod_1608.get(0);
        mod_1609.put(0, t);
    endrule
    rule rule_2076;
        ChannelMessage t;
        t <- mod_1637.get(0);
        mod_1607.put(1, t);
    endrule
    rule rule_2077;
        ChannelMessage t;
        t <- mod_1627.get(0);
        mod_1628.put(0, t);
    endrule
    rule rule_2078;
        ChannelMessage t;
        t <- mod_1638.get(0);
        mod_1605.put(1, t);
    endrule
    rule rule_2079;
        ChannelMessage t;
        t <- mod_1634.get(0);
        mod_1633.put(1, t);
    endrule
    rule rule_2080;
        ChannelMessage t;
        t <- mod_1607.get(1);
        mod_1608.put(0, t);
    endrule
    rule rule_2081;
        ChannelMessage t;
        t <- mod_1619.get(1);
        mod_1612.put(1, t);
    endrule
    rule rule_2082;
        ChannelMessage t;
        t <- mod_1605.get(0);
        mod_1638.put(0, t);
    endrule
    rule rule_2083;
        ChannelMessage t;
        t <- mod_1633.get(1);
        mod_1608.put(1, t);
    endrule
    rule rule_2084;
        ChannelMessage t;
        t <- mod_1635.get(0);
        mod_1633.put(0, t);
    endrule
    rule rule_2085;
        ChannelMessage t;
        t <- mod_1603.get(1);
        mod_1604.put(0, t);
    endrule
    rule rule_2086;
        ChannelMessage t;
        t <- mod_1611.get(1);
        mod_1612.put(0, t);
    endrule
    rule rule_2087;
        ChannelMessage t;
        t <- mod_1620.get(0);
        mod_1619.put(1, t);
    endrule
    rule rule_2088;
        ChannelMessage t;
        t <- mod_1628.get(0);
        mod_1627.put(1, t);
    endrule
    rule rule_2089;
        ChannelMessage t;
        t <- mod_1639.get(1);
        mod_1603.put(1, t);
    endrule
    rule rule_2090;
        ChannelMessage t;
        t <- mod_1639.get(0);
        mod_1639.put(1, t);
    endrule
    rule rule_2091;
        ChannelMessage t;
        t <- mod_1609.get(0);
        mod_1610.put(0, t);
    endrule
    rule rule_2092;
        ChannelMessage t;
        t <- mod_1621.get(0);
        mod_1619.put(0, t);
    endrule
    rule rule_2093;
        ChannelMessage t;
        t <- mod_1605.get(1);
        mod_1606.put(0, t);
    endrule
    rule rule_2094;
        ChannelMessage t;
        t <- mod_1632.get(0);
        mod_1631.put(1, t);
    endrule
    rule rule_2095;
        ChannelMessage t;
        t <- mod_1601.get(0);
        mod_1602.put(0, t);
    endrule
    rule rule_2096;
        ChannelMessage t;
        t <- mod_1614.get(1);
        mod_1615.put(0, t);
    endrule
    rule rule_2097;
        ChannelMessage t;
        t <- mod_1606.get(0);
        mod_1631.put(0, t);
    endrule
    rule rule_2098;
        ChannelMessage t;
        t <- mod_1625.get(0);
        mod_1624.put(0, t);
    endrule
    rule rule_2099;
        ChannelMessage t;
        t <- mod_1630.get(0);
        mod_1629.put(0, t);
    endrule
    rule rule_2100;
        ChannelMessage t;
        t <- mod_1636.get(0);
        mod_1635.put(0, t);
    endrule
    rule rule_2101;
        ChannelMessage t;
        t <- mod_1602.get(0);
        mod_1603.put(0, t);
    endrule
    rule rule_2102;
        ChannelMessage t;
        t <- mod_1624.get(0);
        mod_1610.put(1, t);
    endrule
    rule rule_2103;
        ChannelMessage t;
        t <- mod_1610.get(0);
        mod_1611.put(0, t);
    endrule
    rule rule_2104;
        ChannelMessage t;
        t <- mod_1631.get(1);
        mod_1626.put(0, t);
    endrule
    rule rule_2105;
        ChannelMessage t;
        t <- mod_1627.get(1);
        mod_1626.put(1, t);
    endrule
    rule rule_2106;
        ChannelMessage t;
        t <- mod_1622.get(0);
        mod_1621.put(0, t);
    endrule
    rule rule_2107;
        ChannelMessage t;
        t <- mod_1603.get(0);
        mod_1639.put(0, t);
    endrule
    rule rule_2108;
        ChannelMessage t;
        t <- mod_1615.get(1);
        mod_1616.put(1, t);
    endrule
    rule rule_2109;
        ChannelMessage t;
        t <- mod_1617.get(1);
        mod_1615.put(1, t);
    endrule
    rule rule_2110;
        ChannelMessage t;
        t <- mod_1631.get(0);
        mod_1632.put(0, t);
    endrule
    rule rule_2111;
        ChannelMessage t;
        t <- mod_1604.get(3);
        mod_1605.put(0, t);
    endrule
    rule rule_2112;
        ChannelMessage t;
        t <- mod_1606.get(1);
        mod_1607.put(0, t);
    endrule
    rule rule_2113;
        ChannelMessage t;
        t <- mod_1607.get(0);
        mod_1637.put(0, t);
    endrule
    rule rule_2114;
        ChannelMessage t;
        t <- mod_1600.get(0);
        mod_1601.put(0, t);
    endrule
    rule rule_2115;
        ChannelMessage t;
        t <- mod_1623.get(0);
        mod_1611.put(1, t);
    endrule
    rule rule_2116;
        ChannelMessage t;
        t <- mod_1617.get(0);
        mod_1617.put(1, t);
    endrule
    rule rule_2117;
        ChannelMessage t;
        t <- mod_1633.get(0);
        mod_1634.put(0, t);
    endrule
    rule rule_2118;
        ChannelMessage t;
        t <- mod_1618.get(0);
        mod_1618.put(1, t);
    endrule
    rule rule_2119;
        ChannelMessage t;
        t <- mod_1629.get(0);
        mod_1627.put(0, t);
    endrule
    rule rule_2120;
        ChannelMessage t;
        t <- mod_1626.get(0);
        mod_1625.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1600.put(0, t);
        end
        if (i == 1) begin
            mod_1616.put(0, t);
        end
        if (i == 2) begin
            mod_1622.put(0, t);
        end
        if (i == 3) begin
            mod_1630.put(0, t);
        end
        if (i == 4) begin
            mod_1636.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_1604.get(0);
        end
        if (i == 3) begin
            t <- mod_1604.get(1);
        end
        if (i == 0) begin
            t <- mod_1604.get(2);
        end
        if (i == 2) begin
            t <- mod_1616.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6074 (Operation_IFC);
    Operation_IFC mod_1641_inner <- mkReshape(2, 64);
    Operation_IFC mod_1641 <- mkDebugOperation(mod_1641_inner, "mod_1641");
    Operation_IFC mod_1642_inner <- mkFlatten(1);
    Operation_IFC mod_1642 <- mkDebugOperation(mod_1642_inner, "mod_1642");
    Operation_IFC mod_1643_inner <- mkFlatten(2);
    Operation_IFC mod_1643 <- mkDebugOperation(mod_1643_inner, "mod_1643");
    Operation_IFC mod_1644_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1644 <- mkDebugOperation(mod_1644_inner, "mod_1644");
    Broadcast_IFC#(4) mod_1645_inner <- mkBroadcast(4);
    Operation_IFC mod_1645 <- mkDebugOperation(mod_1645_inner.op, "mod_1645");
    PMU_IFC mod_1646_bufferize <- mkPMU(2);
    Operation_IFC mod_1646_inner = mod_1646_bufferize.operation;
    Operation_IFC mod_1646 <- mkDebugOperation(mod_1646_inner, "mod_1646");
    Broadcast_IFC#(2) mod_1647_inner <- mkBroadcast(2);
    Operation_IFC mod_1647 <- mkDebugOperation(mod_1647_inner.op, "mod_1647");
    PMU_IFC mod_1648_bufferize <- mkPMU(1);
    Operation_IFC mod_1648_inner = mod_1648_bufferize.operation;
    Operation_IFC mod_1648 <- mkDebugOperation(mod_1648_inner, "mod_1648");
    Operation_IFC mod_1649_inner <- mkBinaryMap(1116, matmul_t_tile);
    Operation_IFC mod_1649 <- mkDebugOperation(mod_1649_inner, "mod_1649");
    Operation_IFC mod_1650_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1650 <- mkDebugOperation(mod_1650_inner, "mod_1650");
    Operation_IFC mod_1651_inner <- mkBinaryMap(1884, mul_tile);
    Operation_IFC mod_1651 <- mkDebugOperation(mod_1651_inner, "mod_1651");
    PMU_IFC mod_1652_bufferize <- mkPMU(1);
    Operation_IFC mod_1652_inner = mod_1652_bufferize.operation;
    Operation_IFC mod_1652 <- mkDebugOperation(mod_1652_inner, "mod_1652");
    Operation_IFC mod_1653_inner <- mkBinaryMap(2483, matmul_t_tile);
    Operation_IFC mod_1653 <- mkDebugOperation(mod_1653_inner, "mod_1653");
    Operation_IFC mod_1654_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1654 <- mkDebugOperation(mod_1654_inner, "mod_1654");
    Operation_IFC mod_1655_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1655 <- mkDebugOperation(mod_1655_inner, "mod_1655");
    Operation_IFC mod_1656_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1656 <- mkDebugOperation(mod_1656_inner, "mod_1656");
    Operation_IFC mod_1657_inner <- mkBinaryMap(2783, mul_tile);
    Operation_IFC mod_1657 <- mkDebugOperation(mod_1657_inner, "mod_1657");
    PMU_IFC mod_1658_bufferize <- mkPMU(1);
    Operation_IFC mod_1658_inner = mod_1658_bufferize.operation;
    Operation_IFC mod_1658 <- mkDebugOperation(mod_1658_inner, "mod_1658");
    PMU_IFC mod_1659_bufferize <- mkPMU(2);
    Operation_IFC mod_1659_inner = mod_1659_bufferize.operation;
    Operation_IFC mod_1659 <- mkDebugOperation(mod_1659_inner, "mod_1659");
    PMU_IFC mod_1660_bufferize <- mkPMU(2);
    Operation_IFC mod_1660_inner = mod_1660_bufferize.operation;
    Operation_IFC mod_1660 <- mkDebugOperation(mod_1660_inner, "mod_1660");
    Operation_IFC mod_1661_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1661 <- mkDebugOperation(mod_1661_inner, "mod_1661");
    Operation_IFC mod_1662_inner <- mkFlatten(1);
    Operation_IFC mod_1662 <- mkDebugOperation(mod_1662_inner, "mod_1662");
    Operation_IFC mod_1663_inner <- mkFlatten(0);
    Operation_IFC mod_1663 <- mkDebugOperation(mod_1663_inner, "mod_1663");
    Operation_IFC mod_1664_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1664 <- mkDebugOperation(mod_1664_inner, "mod_1664");
    Operation_IFC mod_1665_inner <- mkUnaryMap(1756, silu_tile);
    Operation_IFC mod_1665 <- mkDebugOperation(mod_1665_inner, "mod_1665");
    Operation_IFC mod_1666_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1666 <- mkDebugOperation(mod_1666_inner, "mod_1666");
    Operation_IFC mod_1667_inner <- mkBinaryMap(1628, matmul_t_tile);
    Operation_IFC mod_1667 <- mkDebugOperation(mod_1667_inner, "mod_1667");
    PMU_IFC mod_1668_bufferize <- mkPMU(2);
    Operation_IFC mod_1668_inner = mod_1668_bufferize.operation;
    Operation_IFC mod_1668 <- mkDebugOperation(mod_1668_inner, "mod_1668");
    Operation_IFC mod_1669_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1669 <- mkDebugOperation(mod_1669_inner, "mod_1669");
    Operation_IFC mod_1670_inner <- mkFlatten(1);
    Operation_IFC mod_1670 <- mkDebugOperation(mod_1670_inner, "mod_1670");
    Operation_IFC mod_1671_inner <- mkFlatten(0);
    Operation_IFC mod_1671 <- mkDebugOperation(mod_1671_inner, "mod_1671");
    PMU_IFC mod_1672_bufferize <- mkPMU(1);
    Operation_IFC mod_1672_inner = mod_1672_bufferize.operation;
    Operation_IFC mod_1672 <- mkDebugOperation(mod_1672_inner, "mod_1672");
    Operation_IFC mod_1673_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1673 <- mkDebugOperation(mod_1673_inner, "mod_1673");
    PMU_IFC mod_1674_bufferize <- mkPMU(2);
    Operation_IFC mod_1674_inner = mod_1674_bufferize.operation;
    Operation_IFC mod_1674 <- mkDebugOperation(mod_1674_inner, "mod_1674");
    Operation_IFC mod_1675_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1675 <- mkDebugOperation(mod_1675_inner, "mod_1675");
    Operation_IFC mod_1676_inner <- mkFlatten(1);
    Operation_IFC mod_1676 <- mkDebugOperation(mod_1676_inner, "mod_1676");
    Operation_IFC mod_1677_inner <- mkFlatten(0);
    Operation_IFC mod_1677 <- mkDebugOperation(mod_1677_inner, "mod_1677");
    Operation_IFC mod_1678_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1678 <- mkDebugOperation(mod_1678_inner, "mod_1678");
    Operation_IFC mod_1679_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1679 <- mkDebugOperation(mod_1679_inner, "mod_1679");
    PMU_IFC mod_1680_bufferize <- mkPMU(2);
    Operation_IFC mod_1680_inner = mod_1680_bufferize.operation;
    Operation_IFC mod_1680 <- mkDebugOperation(mod_1680_inner, "mod_1680");
    rule rule_2121;
        ChannelMessage t;
        t <- mod_1664.get(0);
        mod_1652.put(1, t);
    endrule
    rule rule_2122;
        ChannelMessage t;
        t <- mod_1669.get(0);
        mod_1668.put(1, t);
    endrule
    rule rule_2123;
        ChannelMessage t;
        t <- mod_1648.get(1);
        mod_1649.put(0, t);
    endrule
    rule rule_2124;
        ChannelMessage t;
        t <- mod_1660.get(1);
        mod_1653.put(1, t);
    endrule
    rule rule_2125;
        ChannelMessage t;
        t <- mod_1662.get(0);
        mod_1660.put(0, t);
    endrule
    rule rule_2126;
        ChannelMessage t;
        t <- mod_1670.get(0);
        mod_1668.put(0, t);
    endrule
    rule rule_2127;
        ChannelMessage t;
        t <- mod_1643.get(0);
        mod_1644.put(0, t);
    endrule
    rule rule_2128;
        ChannelMessage t;
        t <- mod_1644.get(0);
        mod_1680.put(0, t);
    endrule
    rule rule_2129;
        ChannelMessage t;
        t <- mod_1673.get(0);
        mod_1672.put(1, t);
    endrule
    rule rule_2130;
        ChannelMessage t;
        t <- mod_1652.get(1);
        mod_1653.put(0, t);
    endrule
    rule rule_2131;
        ChannelMessage t;
        t <- mod_1680.get(0);
        mod_1680.put(1, t);
    endrule
    rule rule_2132;
        ChannelMessage t;
        t <- mod_1642.get(0);
        mod_1643.put(0, t);
    endrule
    rule rule_2133;
        ChannelMessage t;
        t <- mod_1661.get(0);
        mod_1660.put(1, t);
    endrule
    rule rule_2134;
        ChannelMessage t;
        t <- mod_1641.get(0);
        mod_1642.put(0, t);
    endrule
    rule rule_2135;
        ChannelMessage t;
        t <- mod_1676.get(0);
        mod_1674.put(0, t);
    endrule
    rule rule_2136;
        ChannelMessage t;
        t <- mod_1677.get(0);
        mod_1676.put(0, t);
    endrule
    rule rule_2137;
        ChannelMessage t;
        t <- mod_1659.get(0);
        mod_1659.put(1, t);
    endrule
    rule rule_2138;
        ChannelMessage t;
        t <- mod_1659.get(1);
        mod_1655.put(1, t);
    endrule
    rule rule_2139;
        ChannelMessage t;
        t <- mod_1663.get(0);
        mod_1662.put(0, t);
    endrule
    rule rule_2140;
        ChannelMessage t;
        t <- mod_1660.get(0);
        mod_1661.put(0, t);
    endrule
    rule rule_2141;
        ChannelMessage t;
        t <- mod_1652.get(0);
        mod_1664.put(0, t);
    endrule
    rule rule_2142;
        ChannelMessage t;
        t <- mod_1672.get(1);
        mod_1667.put(0, t);
    endrule
    rule rule_2143;
        ChannelMessage t;
        t <- mod_1678.get(0);
        mod_1648.put(1, t);
    endrule
    rule rule_2144;
        ChannelMessage t;
        t <- mod_1651.get(0);
        mod_1652.put(0, t);
    endrule
    rule rule_2145;
        ChannelMessage t;
        t <- mod_1649.get(0);
        mod_1650.put(0, t);
    endrule
    rule rule_2146;
        ChannelMessage t;
        t <- mod_1674.get(0);
        mod_1675.put(0, t);
    endrule
    rule rule_2147;
        ChannelMessage t;
        t <- mod_1666.get(0);
        mod_1665.put(0, t);
    endrule
    rule rule_2148;
        ChannelMessage t;
        t <- mod_1674.get(1);
        mod_1649.put(1, t);
    endrule
    rule rule_2149;
        ChannelMessage t;
        t <- mod_1679.get(0);
        mod_1646.put(1, t);
    endrule
    rule rule_2150;
        ChannelMessage t;
        t <- mod_1658.get(0);
        mod_1658.put(1, t);
    endrule
    rule rule_2151;
        ChannelMessage t;
        t <- mod_1656.get(1);
        mod_1657.put(1, t);
    endrule
    rule rule_2152;
        ChannelMessage t;
        t <- mod_1668.get(1);
        mod_1667.put(1, t);
    endrule
    rule rule_2153;
        ChannelMessage t;
        t <- mod_1646.get(0);
        mod_1679.put(0, t);
    endrule
    rule rule_2154;
        ChannelMessage t;
        t <- mod_1655.get(1);
        mod_1656.put(0, t);
    endrule
    rule rule_2155;
        ChannelMessage t;
        t <- mod_1668.get(0);
        mod_1669.put(0, t);
    endrule
    rule rule_2156;
        ChannelMessage t;
        t <- mod_1646.get(1);
        mod_1647.put(0, t);
    endrule
    rule rule_2157;
        ChannelMessage t;
        t <- mod_1658.get(1);
        mod_1656.put(1, t);
    endrule
    rule rule_2158;
        ChannelMessage t;
        t <- mod_1672.get(0);
        mod_1673.put(0, t);
    endrule
    rule rule_2159;
        ChannelMessage t;
        t <- mod_1644.get(1);
        mod_1645.put(0, t);
    endrule
    rule rule_2160;
        ChannelMessage t;
        t <- mod_1655.get(0);
        mod_1659.put(0, t);
    endrule
    rule rule_2161;
        ChannelMessage t;
        t <- mod_1653.get(0);
        mod_1654.put(0, t);
    endrule
    rule rule_2162;
        ChannelMessage t;
        t <- mod_1675.get(0);
        mod_1674.put(1, t);
    endrule
    rule rule_2163;
        ChannelMessage t;
        t <- mod_1647.get(0);
        mod_1672.put(0, t);
    endrule
    rule rule_2164;
        ChannelMessage t;
        t <- mod_1650.get(0);
        mod_1651.put(0, t);
    endrule
    rule rule_2165;
        ChannelMessage t;
        t <- mod_1667.get(0);
        mod_1666.put(0, t);
    endrule
    rule rule_2166;
        ChannelMessage t;
        t <- mod_1656.get(0);
        mod_1658.put(0, t);
    endrule
    rule rule_2167;
        ChannelMessage t;
        t <- mod_1648.get(0);
        mod_1678.put(0, t);
    endrule
    rule rule_2168;
        ChannelMessage t;
        t <- mod_1671.get(0);
        mod_1670.put(0, t);
    endrule
    rule rule_2169;
        ChannelMessage t;
        t <- mod_1647.get(1);
        mod_1648.put(0, t);
    endrule
    rule rule_2170;
        ChannelMessage t;
        t <- mod_1665.get(0);
        mod_1651.put(1, t);
    endrule
    rule rule_2171;
        ChannelMessage t;
        t <- mod_1645.get(3);
        mod_1646.put(0, t);
    endrule
    rule rule_2172;
        ChannelMessage t;
        t <- mod_1654.get(0);
        mod_1655.put(0, t);
    endrule
    rule rule_2173;
        ChannelMessage t;
        t <- mod_1680.get(1);
        mod_1644.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1641.put(0, t);
        end
        if (i == 1) begin
            mod_1657.put(0, t);
        end
        if (i == 2) begin
            mod_1663.put(0, t);
        end
        if (i == 3) begin
            mod_1671.put(0, t);
        end
        if (i == 4) begin
            mod_1677.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 2) begin
            t <- mod_1645.get(0);
        end
        if (i == 1) begin
            t <- mod_1645.get(1);
        end
        if (i == 0) begin
            t <- mod_1645.get(2);
        end
        if (i == 3) begin
            t <- mod_1657.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6075 (Operation_IFC);
    Operation_IFC mod_1682_inner <- mkReshape(2, 64);
    Operation_IFC mod_1682 <- mkDebugOperation(mod_1682_inner, "mod_1682");
    Operation_IFC mod_1683_inner <- mkFlatten(1);
    Operation_IFC mod_1683 <- mkDebugOperation(mod_1683_inner, "mod_1683");
    Operation_IFC mod_1684_inner <- mkFlatten(2);
    Operation_IFC mod_1684 <- mkDebugOperation(mod_1684_inner, "mod_1684");
    Operation_IFC mod_1685_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1685 <- mkDebugOperation(mod_1685_inner, "mod_1685");
    Broadcast_IFC#(4) mod_1686_inner <- mkBroadcast(4);
    Operation_IFC mod_1686 <- mkDebugOperation(mod_1686_inner.op, "mod_1686");
    PMU_IFC mod_1687_bufferize <- mkPMU(2);
    Operation_IFC mod_1687_inner = mod_1687_bufferize.operation;
    Operation_IFC mod_1687 <- mkDebugOperation(mod_1687_inner, "mod_1687");
    Broadcast_IFC#(2) mod_1688_inner <- mkBroadcast(2);
    Operation_IFC mod_1688 <- mkDebugOperation(mod_1688_inner.op, "mod_1688");
    PMU_IFC mod_1689_bufferize <- mkPMU(1);
    Operation_IFC mod_1689_inner = mod_1689_bufferize.operation;
    Operation_IFC mod_1689 <- mkDebugOperation(mod_1689_inner, "mod_1689");
    Operation_IFC mod_1690_inner <- mkBinaryMap(1115, matmul_t_tile);
    Operation_IFC mod_1690 <- mkDebugOperation(mod_1690_inner, "mod_1690");
    Operation_IFC mod_1691_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1691 <- mkDebugOperation(mod_1691_inner, "mod_1691");
    Operation_IFC mod_1692_inner <- mkBinaryMap(1883, mul_tile);
    Operation_IFC mod_1692 <- mkDebugOperation(mod_1692_inner, "mod_1692");
    PMU_IFC mod_1693_bufferize <- mkPMU(1);
    Operation_IFC mod_1693_inner = mod_1693_bufferize.operation;
    Operation_IFC mod_1693 <- mkDebugOperation(mod_1693_inner, "mod_1693");
    Operation_IFC mod_1694_inner <- mkBinaryMap(2481, matmul_t_tile);
    Operation_IFC mod_1694 <- mkDebugOperation(mod_1694_inner, "mod_1694");
    Operation_IFC mod_1695_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1695 <- mkDebugOperation(mod_1695_inner, "mod_1695");
    Operation_IFC mod_1696_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1696 <- mkDebugOperation(mod_1696_inner, "mod_1696");
    Operation_IFC mod_1697_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1697 <- mkDebugOperation(mod_1697_inner, "mod_1697");
    Operation_IFC mod_1698_inner <- mkBinaryMap(2782, mul_tile);
    Operation_IFC mod_1698 <- mkDebugOperation(mod_1698_inner, "mod_1698");
    PMU_IFC mod_1699_bufferize <- mkPMU(1);
    Operation_IFC mod_1699_inner = mod_1699_bufferize.operation;
    Operation_IFC mod_1699 <- mkDebugOperation(mod_1699_inner, "mod_1699");
    PMU_IFC mod_1700_bufferize <- mkPMU(2);
    Operation_IFC mod_1700_inner = mod_1700_bufferize.operation;
    Operation_IFC mod_1700 <- mkDebugOperation(mod_1700_inner, "mod_1700");
    PMU_IFC mod_1701_bufferize <- mkPMU(2);
    Operation_IFC mod_1701_inner = mod_1701_bufferize.operation;
    Operation_IFC mod_1701 <- mkDebugOperation(mod_1701_inner, "mod_1701");
    Operation_IFC mod_1702_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1702 <- mkDebugOperation(mod_1702_inner, "mod_1702");
    Operation_IFC mod_1703_inner <- mkFlatten(1);
    Operation_IFC mod_1703 <- mkDebugOperation(mod_1703_inner, "mod_1703");
    Operation_IFC mod_1704_inner <- mkFlatten(0);
    Operation_IFC mod_1704 <- mkDebugOperation(mod_1704_inner, "mod_1704");
    Operation_IFC mod_1705_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1705 <- mkDebugOperation(mod_1705_inner, "mod_1705");
    Operation_IFC mod_1706_inner <- mkUnaryMap(1755, silu_tile);
    Operation_IFC mod_1706 <- mkDebugOperation(mod_1706_inner, "mod_1706");
    Operation_IFC mod_1707_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1707 <- mkDebugOperation(mod_1707_inner, "mod_1707");
    Operation_IFC mod_1708_inner <- mkBinaryMap(1627, matmul_t_tile);
    Operation_IFC mod_1708 <- mkDebugOperation(mod_1708_inner, "mod_1708");
    PMU_IFC mod_1709_bufferize <- mkPMU(2);
    Operation_IFC mod_1709_inner = mod_1709_bufferize.operation;
    Operation_IFC mod_1709 <- mkDebugOperation(mod_1709_inner, "mod_1709");
    Operation_IFC mod_1710_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1710 <- mkDebugOperation(mod_1710_inner, "mod_1710");
    Operation_IFC mod_1711_inner <- mkFlatten(1);
    Operation_IFC mod_1711 <- mkDebugOperation(mod_1711_inner, "mod_1711");
    Operation_IFC mod_1712_inner <- mkFlatten(0);
    Operation_IFC mod_1712 <- mkDebugOperation(mod_1712_inner, "mod_1712");
    PMU_IFC mod_1713_bufferize <- mkPMU(1);
    Operation_IFC mod_1713_inner = mod_1713_bufferize.operation;
    Operation_IFC mod_1713 <- mkDebugOperation(mod_1713_inner, "mod_1713");
    Operation_IFC mod_1714_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1714 <- mkDebugOperation(mod_1714_inner, "mod_1714");
    PMU_IFC mod_1715_bufferize <- mkPMU(2);
    Operation_IFC mod_1715_inner = mod_1715_bufferize.operation;
    Operation_IFC mod_1715 <- mkDebugOperation(mod_1715_inner, "mod_1715");
    Operation_IFC mod_1716_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1716 <- mkDebugOperation(mod_1716_inner, "mod_1716");
    Operation_IFC mod_1717_inner <- mkFlatten(1);
    Operation_IFC mod_1717 <- mkDebugOperation(mod_1717_inner, "mod_1717");
    Operation_IFC mod_1718_inner <- mkFlatten(0);
    Operation_IFC mod_1718 <- mkDebugOperation(mod_1718_inner, "mod_1718");
    Operation_IFC mod_1719_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1719 <- mkDebugOperation(mod_1719_inner, "mod_1719");
    Operation_IFC mod_1720_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1720 <- mkDebugOperation(mod_1720_inner, "mod_1720");
    PMU_IFC mod_1721_bufferize <- mkPMU(2);
    Operation_IFC mod_1721_inner = mod_1721_bufferize.operation;
    Operation_IFC mod_1721 <- mkDebugOperation(mod_1721_inner, "mod_1721");
    rule rule_2174;
        ChannelMessage t;
        t <- mod_1688.get(1);
        mod_1689.put(0, t);
    endrule
    rule rule_2175;
        ChannelMessage t;
        t <- mod_1697.get(0);
        mod_1699.put(0, t);
    endrule
    rule rule_2176;
        ChannelMessage t;
        t <- mod_1682.get(0);
        mod_1683.put(0, t);
    endrule
    rule rule_2177;
        ChannelMessage t;
        t <- mod_1696.get(1);
        mod_1697.put(0, t);
    endrule
    rule rule_2178;
        ChannelMessage t;
        t <- mod_1702.get(0);
        mod_1701.put(1, t);
    endrule
    rule rule_2179;
        ChannelMessage t;
        t <- mod_1711.get(0);
        mod_1709.put(0, t);
    endrule
    rule rule_2180;
        ChannelMessage t;
        t <- mod_1706.get(0);
        mod_1692.put(1, t);
    endrule
    rule rule_2181;
        ChannelMessage t;
        t <- mod_1699.get(1);
        mod_1697.put(1, t);
    endrule
    rule rule_2182;
        ChannelMessage t;
        t <- mod_1704.get(0);
        mod_1703.put(0, t);
    endrule
    rule rule_2183;
        ChannelMessage t;
        t <- mod_1687.get(1);
        mod_1688.put(0, t);
    endrule
    rule rule_2184;
        ChannelMessage t;
        t <- mod_1685.get(0);
        mod_1721.put(0, t);
    endrule
    rule rule_2185;
        ChannelMessage t;
        t <- mod_1685.get(1);
        mod_1686.put(0, t);
    endrule
    rule rule_2186;
        ChannelMessage t;
        t <- mod_1695.get(0);
        mod_1696.put(0, t);
    endrule
    rule rule_2187;
        ChannelMessage t;
        t <- mod_1716.get(0);
        mod_1715.put(1, t);
    endrule
    rule rule_2188;
        ChannelMessage t;
        t <- mod_1689.get(0);
        mod_1719.put(0, t);
    endrule
    rule rule_2189;
        ChannelMessage t;
        t <- mod_1703.get(0);
        mod_1701.put(0, t);
    endrule
    rule rule_2190;
        ChannelMessage t;
        t <- mod_1690.get(0);
        mod_1691.put(0, t);
    endrule
    rule rule_2191;
        ChannelMessage t;
        t <- mod_1718.get(0);
        mod_1717.put(0, t);
    endrule
    rule rule_2192;
        ChannelMessage t;
        t <- mod_1696.get(0);
        mod_1700.put(0, t);
    endrule
    rule rule_2193;
        ChannelMessage t;
        t <- mod_1717.get(0);
        mod_1715.put(0, t);
    endrule
    rule rule_2194;
        ChannelMessage t;
        t <- mod_1686.get(3);
        mod_1687.put(0, t);
    endrule
    rule rule_2195;
        ChannelMessage t;
        t <- mod_1709.get(1);
        mod_1708.put(1, t);
    endrule
    rule rule_2196;
        ChannelMessage t;
        t <- mod_1687.get(0);
        mod_1720.put(0, t);
    endrule
    rule rule_2197;
        ChannelMessage t;
        t <- mod_1714.get(0);
        mod_1713.put(1, t);
    endrule
    rule rule_2198;
        ChannelMessage t;
        t <- mod_1709.get(0);
        mod_1710.put(0, t);
    endrule
    rule rule_2199;
        ChannelMessage t;
        t <- mod_1715.get(0);
        mod_1716.put(0, t);
    endrule
    rule rule_2200;
        ChannelMessage t;
        t <- mod_1710.get(0);
        mod_1709.put(1, t);
    endrule
    rule rule_2201;
        ChannelMessage t;
        t <- mod_1721.get(0);
        mod_1721.put(1, t);
    endrule
    rule rule_2202;
        ChannelMessage t;
        t <- mod_1701.get(1);
        mod_1694.put(1, t);
    endrule
    rule rule_2203;
        ChannelMessage t;
        t <- mod_1699.get(0);
        mod_1699.put(1, t);
    endrule
    rule rule_2204;
        ChannelMessage t;
        t <- mod_1692.get(0);
        mod_1693.put(0, t);
    endrule
    rule rule_2205;
        ChannelMessage t;
        t <- mod_1713.get(1);
        mod_1708.put(0, t);
    endrule
    rule rule_2206;
        ChannelMessage t;
        t <- mod_1693.get(1);
        mod_1694.put(0, t);
    endrule
    rule rule_2207;
        ChannelMessage t;
        t <- mod_1693.get(0);
        mod_1705.put(0, t);
    endrule
    rule rule_2208;
        ChannelMessage t;
        t <- mod_1688.get(0);
        mod_1713.put(0, t);
    endrule
    rule rule_2209;
        ChannelMessage t;
        t <- mod_1713.get(0);
        mod_1714.put(0, t);
    endrule
    rule rule_2210;
        ChannelMessage t;
        t <- mod_1715.get(1);
        mod_1690.put(1, t);
    endrule
    rule rule_2211;
        ChannelMessage t;
        t <- mod_1700.get(0);
        mod_1700.put(1, t);
    endrule
    rule rule_2212;
        ChannelMessage t;
        t <- mod_1705.get(0);
        mod_1693.put(1, t);
    endrule
    rule rule_2213;
        ChannelMessage t;
        t <- mod_1691.get(0);
        mod_1692.put(0, t);
    endrule
    rule rule_2214;
        ChannelMessage t;
        t <- mod_1694.get(0);
        mod_1695.put(0, t);
    endrule
    rule rule_2215;
        ChannelMessage t;
        t <- mod_1683.get(0);
        mod_1684.put(0, t);
    endrule
    rule rule_2216;
        ChannelMessage t;
        t <- mod_1701.get(0);
        mod_1702.put(0, t);
    endrule
    rule rule_2217;
        ChannelMessage t;
        t <- mod_1697.get(1);
        mod_1698.put(1, t);
    endrule
    rule rule_2218;
        ChannelMessage t;
        t <- mod_1707.get(0);
        mod_1706.put(0, t);
    endrule
    rule rule_2219;
        ChannelMessage t;
        t <- mod_1708.get(0);
        mod_1707.put(0, t);
    endrule
    rule rule_2220;
        ChannelMessage t;
        t <- mod_1700.get(1);
        mod_1696.put(1, t);
    endrule
    rule rule_2221;
        ChannelMessage t;
        t <- mod_1721.get(1);
        mod_1685.put(1, t);
    endrule
    rule rule_2222;
        ChannelMessage t;
        t <- mod_1712.get(0);
        mod_1711.put(0, t);
    endrule
    rule rule_2223;
        ChannelMessage t;
        t <- mod_1689.get(1);
        mod_1690.put(0, t);
    endrule
    rule rule_2224;
        ChannelMessage t;
        t <- mod_1720.get(0);
        mod_1687.put(1, t);
    endrule
    rule rule_2225;
        ChannelMessage t;
        t <- mod_1684.get(0);
        mod_1685.put(0, t);
    endrule
    rule rule_2226;
        ChannelMessage t;
        t <- mod_1719.get(0);
        mod_1689.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1682.put(0, t);
        end
        if (i == 1) begin
            mod_1698.put(0, t);
        end
        if (i == 2) begin
            mod_1704.put(0, t);
        end
        if (i == 3) begin
            mod_1712.put(0, t);
        end
        if (i == 4) begin
            mod_1718.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_1686.get(0);
        end
        if (i == 0) begin
            t <- mod_1686.get(1);
        end
        if (i == 2) begin
            t <- mod_1686.get(2);
        end
        if (i == 3) begin
            t <- mod_1698.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6076 (Operation_IFC);
    Operation_IFC mod_1723_inner <- mkReshape(2, 64);
    Operation_IFC mod_1723 <- mkDebugOperation(mod_1723_inner, "mod_1723");
    Operation_IFC mod_1724_inner <- mkFlatten(1);
    Operation_IFC mod_1724 <- mkDebugOperation(mod_1724_inner, "mod_1724");
    Operation_IFC mod_1725_inner <- mkFlatten(2);
    Operation_IFC mod_1725 <- mkDebugOperation(mod_1725_inner, "mod_1725");
    Operation_IFC mod_1726_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1726 <- mkDebugOperation(mod_1726_inner, "mod_1726");
    Broadcast_IFC#(4) mod_1727_inner <- mkBroadcast(4);
    Operation_IFC mod_1727 <- mkDebugOperation(mod_1727_inner.op, "mod_1727");
    PMU_IFC mod_1728_bufferize <- mkPMU(2);
    Operation_IFC mod_1728_inner = mod_1728_bufferize.operation;
    Operation_IFC mod_1728 <- mkDebugOperation(mod_1728_inner, "mod_1728");
    Broadcast_IFC#(2) mod_1729_inner <- mkBroadcast(2);
    Operation_IFC mod_1729 <- mkDebugOperation(mod_1729_inner.op, "mod_1729");
    PMU_IFC mod_1730_bufferize <- mkPMU(1);
    Operation_IFC mod_1730_inner = mod_1730_bufferize.operation;
    Operation_IFC mod_1730 <- mkDebugOperation(mod_1730_inner, "mod_1730");
    Operation_IFC mod_1731_inner <- mkBinaryMap(1114, matmul_t_tile);
    Operation_IFC mod_1731 <- mkDebugOperation(mod_1731_inner, "mod_1731");
    Operation_IFC mod_1732_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1732 <- mkDebugOperation(mod_1732_inner, "mod_1732");
    Operation_IFC mod_1733_inner <- mkBinaryMap(1882, mul_tile);
    Operation_IFC mod_1733 <- mkDebugOperation(mod_1733_inner, "mod_1733");
    PMU_IFC mod_1734_bufferize <- mkPMU(1);
    Operation_IFC mod_1734_inner = mod_1734_bufferize.operation;
    Operation_IFC mod_1734 <- mkDebugOperation(mod_1734_inner, "mod_1734");
    Operation_IFC mod_1735_inner <- mkBinaryMap(2479, matmul_t_tile);
    Operation_IFC mod_1735 <- mkDebugOperation(mod_1735_inner, "mod_1735");
    Operation_IFC mod_1736_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1736 <- mkDebugOperation(mod_1736_inner, "mod_1736");
    Operation_IFC mod_1737_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1737 <- mkDebugOperation(mod_1737_inner, "mod_1737");
    Operation_IFC mod_1738_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1738 <- mkDebugOperation(mod_1738_inner, "mod_1738");
    Operation_IFC mod_1739_inner <- mkBinaryMap(2781, mul_tile);
    Operation_IFC mod_1739 <- mkDebugOperation(mod_1739_inner, "mod_1739");
    PMU_IFC mod_1740_bufferize <- mkPMU(1);
    Operation_IFC mod_1740_inner = mod_1740_bufferize.operation;
    Operation_IFC mod_1740 <- mkDebugOperation(mod_1740_inner, "mod_1740");
    PMU_IFC mod_1741_bufferize <- mkPMU(2);
    Operation_IFC mod_1741_inner = mod_1741_bufferize.operation;
    Operation_IFC mod_1741 <- mkDebugOperation(mod_1741_inner, "mod_1741");
    PMU_IFC mod_1742_bufferize <- mkPMU(2);
    Operation_IFC mod_1742_inner = mod_1742_bufferize.operation;
    Operation_IFC mod_1742 <- mkDebugOperation(mod_1742_inner, "mod_1742");
    Operation_IFC mod_1743_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1743 <- mkDebugOperation(mod_1743_inner, "mod_1743");
    Operation_IFC mod_1744_inner <- mkFlatten(1);
    Operation_IFC mod_1744 <- mkDebugOperation(mod_1744_inner, "mod_1744");
    Operation_IFC mod_1745_inner <- mkFlatten(0);
    Operation_IFC mod_1745 <- mkDebugOperation(mod_1745_inner, "mod_1745");
    Operation_IFC mod_1746_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1746 <- mkDebugOperation(mod_1746_inner, "mod_1746");
    Operation_IFC mod_1747_inner <- mkUnaryMap(1754, silu_tile);
    Operation_IFC mod_1747 <- mkDebugOperation(mod_1747_inner, "mod_1747");
    Operation_IFC mod_1748_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1748 <- mkDebugOperation(mod_1748_inner, "mod_1748");
    Operation_IFC mod_1749_inner <- mkBinaryMap(1626, matmul_t_tile);
    Operation_IFC mod_1749 <- mkDebugOperation(mod_1749_inner, "mod_1749");
    PMU_IFC mod_1750_bufferize <- mkPMU(2);
    Operation_IFC mod_1750_inner = mod_1750_bufferize.operation;
    Operation_IFC mod_1750 <- mkDebugOperation(mod_1750_inner, "mod_1750");
    Operation_IFC mod_1751_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1751 <- mkDebugOperation(mod_1751_inner, "mod_1751");
    Operation_IFC mod_1752_inner <- mkFlatten(1);
    Operation_IFC mod_1752 <- mkDebugOperation(mod_1752_inner, "mod_1752");
    Operation_IFC mod_1753_inner <- mkFlatten(0);
    Operation_IFC mod_1753 <- mkDebugOperation(mod_1753_inner, "mod_1753");
    PMU_IFC mod_1754_bufferize <- mkPMU(1);
    Operation_IFC mod_1754_inner = mod_1754_bufferize.operation;
    Operation_IFC mod_1754 <- mkDebugOperation(mod_1754_inner, "mod_1754");
    Operation_IFC mod_1755_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1755 <- mkDebugOperation(mod_1755_inner, "mod_1755");
    PMU_IFC mod_1756_bufferize <- mkPMU(2);
    Operation_IFC mod_1756_inner = mod_1756_bufferize.operation;
    Operation_IFC mod_1756 <- mkDebugOperation(mod_1756_inner, "mod_1756");
    Operation_IFC mod_1757_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1757 <- mkDebugOperation(mod_1757_inner, "mod_1757");
    Operation_IFC mod_1758_inner <- mkFlatten(1);
    Operation_IFC mod_1758 <- mkDebugOperation(mod_1758_inner, "mod_1758");
    Operation_IFC mod_1759_inner <- mkFlatten(0);
    Operation_IFC mod_1759 <- mkDebugOperation(mod_1759_inner, "mod_1759");
    Operation_IFC mod_1760_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1760 <- mkDebugOperation(mod_1760_inner, "mod_1760");
    Operation_IFC mod_1761_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1761 <- mkDebugOperation(mod_1761_inner, "mod_1761");
    PMU_IFC mod_1762_bufferize <- mkPMU(2);
    Operation_IFC mod_1762_inner = mod_1762_bufferize.operation;
    Operation_IFC mod_1762 <- mkDebugOperation(mod_1762_inner, "mod_1762");
    rule rule_2227;
        ChannelMessage t;
        t <- mod_1735.get(0);
        mod_1736.put(0, t);
    endrule
    rule rule_2228;
        ChannelMessage t;
        t <- mod_1746.get(0);
        mod_1734.put(1, t);
    endrule
    rule rule_2229;
        ChannelMessage t;
        t <- mod_1724.get(0);
        mod_1725.put(0, t);
    endrule
    rule rule_2230;
        ChannelMessage t;
        t <- mod_1729.get(0);
        mod_1754.put(0, t);
    endrule
    rule rule_2231;
        ChannelMessage t;
        t <- mod_1728.get(1);
        mod_1729.put(0, t);
    endrule
    rule rule_2232;
        ChannelMessage t;
        t <- mod_1740.get(0);
        mod_1740.put(1, t);
    endrule
    rule rule_2233;
        ChannelMessage t;
        t <- mod_1731.get(0);
        mod_1732.put(0, t);
    endrule
    rule rule_2234;
        ChannelMessage t;
        t <- mod_1742.get(1);
        mod_1735.put(1, t);
    endrule
    rule rule_2235;
        ChannelMessage t;
        t <- mod_1750.get(1);
        mod_1749.put(1, t);
    endrule
    rule rule_2236;
        ChannelMessage t;
        t <- mod_1759.get(0);
        mod_1758.put(0, t);
    endrule
    rule rule_2237;
        ChannelMessage t;
        t <- mod_1758.get(0);
        mod_1756.put(0, t);
    endrule
    rule rule_2238;
        ChannelMessage t;
        t <- mod_1730.get(0);
        mod_1760.put(0, t);
    endrule
    rule rule_2239;
        ChannelMessage t;
        t <- mod_1738.get(1);
        mod_1739.put(1, t);
    endrule
    rule rule_2240;
        ChannelMessage t;
        t <- mod_1723.get(0);
        mod_1724.put(0, t);
    endrule
    rule rule_2241;
        ChannelMessage t;
        t <- mod_1752.get(0);
        mod_1750.put(0, t);
    endrule
    rule rule_2242;
        ChannelMessage t;
        t <- mod_1754.get(0);
        mod_1755.put(0, t);
    endrule
    rule rule_2243;
        ChannelMessage t;
        t <- mod_1756.get(0);
        mod_1757.put(0, t);
    endrule
    rule rule_2244;
        ChannelMessage t;
        t <- mod_1740.get(1);
        mod_1738.put(1, t);
    endrule
    rule rule_2245;
        ChannelMessage t;
        t <- mod_1761.get(0);
        mod_1728.put(1, t);
    endrule
    rule rule_2246;
        ChannelMessage t;
        t <- mod_1754.get(1);
        mod_1749.put(0, t);
    endrule
    rule rule_2247;
        ChannelMessage t;
        t <- mod_1729.get(1);
        mod_1730.put(0, t);
    endrule
    rule rule_2248;
        ChannelMessage t;
        t <- mod_1734.get(0);
        mod_1746.put(0, t);
    endrule
    rule rule_2249;
        ChannelMessage t;
        t <- mod_1732.get(0);
        mod_1733.put(0, t);
    endrule
    rule rule_2250;
        ChannelMessage t;
        t <- mod_1726.get(0);
        mod_1762.put(0, t);
    endrule
    rule rule_2251;
        ChannelMessage t;
        t <- mod_1733.get(0);
        mod_1734.put(0, t);
    endrule
    rule rule_2252;
        ChannelMessage t;
        t <- mod_1734.get(1);
        mod_1735.put(0, t);
    endrule
    rule rule_2253;
        ChannelMessage t;
        t <- mod_1737.get(0);
        mod_1741.put(0, t);
    endrule
    rule rule_2254;
        ChannelMessage t;
        t <- mod_1760.get(0);
        mod_1730.put(1, t);
    endrule
    rule rule_2255;
        ChannelMessage t;
        t <- mod_1736.get(0);
        mod_1737.put(0, t);
    endrule
    rule rule_2256;
        ChannelMessage t;
        t <- mod_1751.get(0);
        mod_1750.put(1, t);
    endrule
    rule rule_2257;
        ChannelMessage t;
        t <- mod_1737.get(1);
        mod_1738.put(0, t);
    endrule
    rule rule_2258;
        ChannelMessage t;
        t <- mod_1757.get(0);
        mod_1756.put(1, t);
    endrule
    rule rule_2259;
        ChannelMessage t;
        t <- mod_1756.get(1);
        mod_1731.put(1, t);
    endrule
    rule rule_2260;
        ChannelMessage t;
        t <- mod_1747.get(0);
        mod_1733.put(1, t);
    endrule
    rule rule_2261;
        ChannelMessage t;
        t <- mod_1748.get(0);
        mod_1747.put(0, t);
    endrule
    rule rule_2262;
        ChannelMessage t;
        t <- mod_1762.get(1);
        mod_1726.put(1, t);
    endrule
    rule rule_2263;
        ChannelMessage t;
        t <- mod_1743.get(0);
        mod_1742.put(1, t);
    endrule
    rule rule_2264;
        ChannelMessage t;
        t <- mod_1744.get(0);
        mod_1742.put(0, t);
    endrule
    rule rule_2265;
        ChannelMessage t;
        t <- mod_1749.get(0);
        mod_1748.put(0, t);
    endrule
    rule rule_2266;
        ChannelMessage t;
        t <- mod_1741.get(0);
        mod_1741.put(1, t);
    endrule
    rule rule_2267;
        ChannelMessage t;
        t <- mod_1745.get(0);
        mod_1744.put(0, t);
    endrule
    rule rule_2268;
        ChannelMessage t;
        t <- mod_1725.get(0);
        mod_1726.put(0, t);
    endrule
    rule rule_2269;
        ChannelMessage t;
        t <- mod_1738.get(0);
        mod_1740.put(0, t);
    endrule
    rule rule_2270;
        ChannelMessage t;
        t <- mod_1762.get(0);
        mod_1762.put(1, t);
    endrule
    rule rule_2271;
        ChannelMessage t;
        t <- mod_1730.get(1);
        mod_1731.put(0, t);
    endrule
    rule rule_2272;
        ChannelMessage t;
        t <- mod_1727.get(3);
        mod_1728.put(0, t);
    endrule
    rule rule_2273;
        ChannelMessage t;
        t <- mod_1728.get(0);
        mod_1761.put(0, t);
    endrule
    rule rule_2274;
        ChannelMessage t;
        t <- mod_1750.get(0);
        mod_1751.put(0, t);
    endrule
    rule rule_2275;
        ChannelMessage t;
        t <- mod_1755.get(0);
        mod_1754.put(1, t);
    endrule
    rule rule_2276;
        ChannelMessage t;
        t <- mod_1742.get(0);
        mod_1743.put(0, t);
    endrule
    rule rule_2277;
        ChannelMessage t;
        t <- mod_1753.get(0);
        mod_1752.put(0, t);
    endrule
    rule rule_2278;
        ChannelMessage t;
        t <- mod_1726.get(1);
        mod_1727.put(0, t);
    endrule
    rule rule_2279;
        ChannelMessage t;
        t <- mod_1741.get(1);
        mod_1737.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1723.put(0, t);
        end
        if (i == 1) begin
            mod_1739.put(0, t);
        end
        if (i == 2) begin
            mod_1745.put(0, t);
        end
        if (i == 3) begin
            mod_1753.put(0, t);
        end
        if (i == 4) begin
            mod_1759.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_1727.get(0);
        end
        if (i == 1) begin
            t <- mod_1727.get(1);
        end
        if (i == 2) begin
            t <- mod_1727.get(2);
        end
        if (i == 0) begin
            t <- mod_1739.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6077 (Operation_IFC);
    Operation_IFC mod_1764_inner <- mkReshape(2, 64);
    Operation_IFC mod_1764 <- mkDebugOperation(mod_1764_inner, "mod_1764");
    Operation_IFC mod_1765_inner <- mkFlatten(1);
    Operation_IFC mod_1765 <- mkDebugOperation(mod_1765_inner, "mod_1765");
    Operation_IFC mod_1766_inner <- mkFlatten(2);
    Operation_IFC mod_1766 <- mkDebugOperation(mod_1766_inner, "mod_1766");
    Operation_IFC mod_1767_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1767 <- mkDebugOperation(mod_1767_inner, "mod_1767");
    Broadcast_IFC#(4) mod_1768_inner <- mkBroadcast(4);
    Operation_IFC mod_1768 <- mkDebugOperation(mod_1768_inner.op, "mod_1768");
    PMU_IFC mod_1769_bufferize <- mkPMU(2);
    Operation_IFC mod_1769_inner = mod_1769_bufferize.operation;
    Operation_IFC mod_1769 <- mkDebugOperation(mod_1769_inner, "mod_1769");
    Broadcast_IFC#(2) mod_1770_inner <- mkBroadcast(2);
    Operation_IFC mod_1770 <- mkDebugOperation(mod_1770_inner.op, "mod_1770");
    PMU_IFC mod_1771_bufferize <- mkPMU(1);
    Operation_IFC mod_1771_inner = mod_1771_bufferize.operation;
    Operation_IFC mod_1771 <- mkDebugOperation(mod_1771_inner, "mod_1771");
    Operation_IFC mod_1772_inner <- mkBinaryMap(1113, matmul_t_tile);
    Operation_IFC mod_1772 <- mkDebugOperation(mod_1772_inner, "mod_1772");
    Operation_IFC mod_1773_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1773 <- mkDebugOperation(mod_1773_inner, "mod_1773");
    Operation_IFC mod_1774_inner <- mkBinaryMap(1881, mul_tile);
    Operation_IFC mod_1774 <- mkDebugOperation(mod_1774_inner, "mod_1774");
    PMU_IFC mod_1775_bufferize <- mkPMU(1);
    Operation_IFC mod_1775_inner = mod_1775_bufferize.operation;
    Operation_IFC mod_1775 <- mkDebugOperation(mod_1775_inner, "mod_1775");
    Operation_IFC mod_1776_inner <- mkBinaryMap(2477, matmul_t_tile);
    Operation_IFC mod_1776 <- mkDebugOperation(mod_1776_inner, "mod_1776");
    Operation_IFC mod_1777_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1777 <- mkDebugOperation(mod_1777_inner, "mod_1777");
    Operation_IFC mod_1778_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1778 <- mkDebugOperation(mod_1778_inner, "mod_1778");
    Operation_IFC mod_1779_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1779 <- mkDebugOperation(mod_1779_inner, "mod_1779");
    Operation_IFC mod_1780_inner <- mkBinaryMap(2780, mul_tile);
    Operation_IFC mod_1780 <- mkDebugOperation(mod_1780_inner, "mod_1780");
    PMU_IFC mod_1781_bufferize <- mkPMU(1);
    Operation_IFC mod_1781_inner = mod_1781_bufferize.operation;
    Operation_IFC mod_1781 <- mkDebugOperation(mod_1781_inner, "mod_1781");
    PMU_IFC mod_1782_bufferize <- mkPMU(2);
    Operation_IFC mod_1782_inner = mod_1782_bufferize.operation;
    Operation_IFC mod_1782 <- mkDebugOperation(mod_1782_inner, "mod_1782");
    PMU_IFC mod_1783_bufferize <- mkPMU(2);
    Operation_IFC mod_1783_inner = mod_1783_bufferize.operation;
    Operation_IFC mod_1783 <- mkDebugOperation(mod_1783_inner, "mod_1783");
    Operation_IFC mod_1784_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1784 <- mkDebugOperation(mod_1784_inner, "mod_1784");
    Operation_IFC mod_1785_inner <- mkFlatten(1);
    Operation_IFC mod_1785 <- mkDebugOperation(mod_1785_inner, "mod_1785");
    Operation_IFC mod_1786_inner <- mkFlatten(0);
    Operation_IFC mod_1786 <- mkDebugOperation(mod_1786_inner, "mod_1786");
    Operation_IFC mod_1787_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1787 <- mkDebugOperation(mod_1787_inner, "mod_1787");
    Operation_IFC mod_1788_inner <- mkUnaryMap(1753, silu_tile);
    Operation_IFC mod_1788 <- mkDebugOperation(mod_1788_inner, "mod_1788");
    Operation_IFC mod_1789_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1789 <- mkDebugOperation(mod_1789_inner, "mod_1789");
    Operation_IFC mod_1790_inner <- mkBinaryMap(1625, matmul_t_tile);
    Operation_IFC mod_1790 <- mkDebugOperation(mod_1790_inner, "mod_1790");
    PMU_IFC mod_1791_bufferize <- mkPMU(2);
    Operation_IFC mod_1791_inner = mod_1791_bufferize.operation;
    Operation_IFC mod_1791 <- mkDebugOperation(mod_1791_inner, "mod_1791");
    Operation_IFC mod_1792_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1792 <- mkDebugOperation(mod_1792_inner, "mod_1792");
    Operation_IFC mod_1793_inner <- mkFlatten(1);
    Operation_IFC mod_1793 <- mkDebugOperation(mod_1793_inner, "mod_1793");
    Operation_IFC mod_1794_inner <- mkFlatten(0);
    Operation_IFC mod_1794 <- mkDebugOperation(mod_1794_inner, "mod_1794");
    PMU_IFC mod_1795_bufferize <- mkPMU(1);
    Operation_IFC mod_1795_inner = mod_1795_bufferize.operation;
    Operation_IFC mod_1795 <- mkDebugOperation(mod_1795_inner, "mod_1795");
    Operation_IFC mod_1796_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1796 <- mkDebugOperation(mod_1796_inner, "mod_1796");
    PMU_IFC mod_1797_bufferize <- mkPMU(2);
    Operation_IFC mod_1797_inner = mod_1797_bufferize.operation;
    Operation_IFC mod_1797 <- mkDebugOperation(mod_1797_inner, "mod_1797");
    Operation_IFC mod_1798_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1798 <- mkDebugOperation(mod_1798_inner, "mod_1798");
    Operation_IFC mod_1799_inner <- mkFlatten(1);
    Operation_IFC mod_1799 <- mkDebugOperation(mod_1799_inner, "mod_1799");
    Operation_IFC mod_1800_inner <- mkFlatten(0);
    Operation_IFC mod_1800 <- mkDebugOperation(mod_1800_inner, "mod_1800");
    Operation_IFC mod_1801_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1801 <- mkDebugOperation(mod_1801_inner, "mod_1801");
    Operation_IFC mod_1802_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1802 <- mkDebugOperation(mod_1802_inner, "mod_1802");
    PMU_IFC mod_1803_bufferize <- mkPMU(2);
    Operation_IFC mod_1803_inner = mod_1803_bufferize.operation;
    Operation_IFC mod_1803 <- mkDebugOperation(mod_1803_inner, "mod_1803");
    rule rule_2280;
        ChannelMessage t;
        t <- mod_1800.get(0);
        mod_1799.put(0, t);
    endrule
    rule rule_2281;
        ChannelMessage t;
        t <- mod_1778.get(1);
        mod_1779.put(0, t);
    endrule
    rule rule_2282;
        ChannelMessage t;
        t <- mod_1803.get(0);
        mod_1803.put(1, t);
    endrule
    rule rule_2283;
        ChannelMessage t;
        t <- mod_1787.get(0);
        mod_1775.put(1, t);
    endrule
    rule rule_2284;
        ChannelMessage t;
        t <- mod_1789.get(0);
        mod_1788.put(0, t);
    endrule
    rule rule_2285;
        ChannelMessage t;
        t <- mod_1799.get(0);
        mod_1797.put(0, t);
    endrule
    rule rule_2286;
        ChannelMessage t;
        t <- mod_1801.get(0);
        mod_1771.put(1, t);
    endrule
    rule rule_2287;
        ChannelMessage t;
        t <- mod_1769.get(0);
        mod_1802.put(0, t);
    endrule
    rule rule_2288;
        ChannelMessage t;
        t <- mod_1798.get(0);
        mod_1797.put(1, t);
    endrule
    rule rule_2289;
        ChannelMessage t;
        t <- mod_1791.get(0);
        mod_1792.put(0, t);
    endrule
    rule rule_2290;
        ChannelMessage t;
        t <- mod_1767.get(0);
        mod_1803.put(0, t);
    endrule
    rule rule_2291;
        ChannelMessage t;
        t <- mod_1765.get(0);
        mod_1766.put(0, t);
    endrule
    rule rule_2292;
        ChannelMessage t;
        t <- mod_1786.get(0);
        mod_1785.put(0, t);
    endrule
    rule rule_2293;
        ChannelMessage t;
        t <- mod_1772.get(0);
        mod_1773.put(0, t);
    endrule
    rule rule_2294;
        ChannelMessage t;
        t <- mod_1794.get(0);
        mod_1793.put(0, t);
    endrule
    rule rule_2295;
        ChannelMessage t;
        t <- mod_1769.get(1);
        mod_1770.put(0, t);
    endrule
    rule rule_2296;
        ChannelMessage t;
        t <- mod_1768.get(3);
        mod_1769.put(0, t);
    endrule
    rule rule_2297;
        ChannelMessage t;
        t <- mod_1771.get(1);
        mod_1772.put(0, t);
    endrule
    rule rule_2298;
        ChannelMessage t;
        t <- mod_1773.get(0);
        mod_1774.put(0, t);
    endrule
    rule rule_2299;
        ChannelMessage t;
        t <- mod_1776.get(0);
        mod_1777.put(0, t);
    endrule
    rule rule_2300;
        ChannelMessage t;
        t <- mod_1781.get(0);
        mod_1781.put(1, t);
    endrule
    rule rule_2301;
        ChannelMessage t;
        t <- mod_1781.get(1);
        mod_1779.put(1, t);
    endrule
    rule rule_2302;
        ChannelMessage t;
        t <- mod_1774.get(0);
        mod_1775.put(0, t);
    endrule
    rule rule_2303;
        ChannelMessage t;
        t <- mod_1775.get(0);
        mod_1787.put(0, t);
    endrule
    rule rule_2304;
        ChannelMessage t;
        t <- mod_1777.get(0);
        mod_1778.put(0, t);
    endrule
    rule rule_2305;
        ChannelMessage t;
        t <- mod_1793.get(0);
        mod_1791.put(0, t);
    endrule
    rule rule_2306;
        ChannelMessage t;
        t <- mod_1795.get(0);
        mod_1796.put(0, t);
    endrule
    rule rule_2307;
        ChannelMessage t;
        t <- mod_1796.get(0);
        mod_1795.put(1, t);
    endrule
    rule rule_2308;
        ChannelMessage t;
        t <- mod_1797.get(1);
        mod_1772.put(1, t);
    endrule
    rule rule_2309;
        ChannelMessage t;
        t <- mod_1788.get(0);
        mod_1774.put(1, t);
    endrule
    rule rule_2310;
        ChannelMessage t;
        t <- mod_1764.get(0);
        mod_1765.put(0, t);
    endrule
    rule rule_2311;
        ChannelMessage t;
        t <- mod_1791.get(1);
        mod_1790.put(1, t);
    endrule
    rule rule_2312;
        ChannelMessage t;
        t <- mod_1792.get(0);
        mod_1791.put(1, t);
    endrule
    rule rule_2313;
        ChannelMessage t;
        t <- mod_1779.get(1);
        mod_1780.put(1, t);
    endrule
    rule rule_2314;
        ChannelMessage t;
        t <- mod_1782.get(0);
        mod_1782.put(1, t);
    endrule
    rule rule_2315;
        ChannelMessage t;
        t <- mod_1783.get(1);
        mod_1776.put(1, t);
    endrule
    rule rule_2316;
        ChannelMessage t;
        t <- mod_1795.get(1);
        mod_1790.put(0, t);
    endrule
    rule rule_2317;
        ChannelMessage t;
        t <- mod_1797.get(0);
        mod_1798.put(0, t);
    endrule
    rule rule_2318;
        ChannelMessage t;
        t <- mod_1771.get(0);
        mod_1801.put(0, t);
    endrule
    rule rule_2319;
        ChannelMessage t;
        t <- mod_1767.get(1);
        mod_1768.put(0, t);
    endrule
    rule rule_2320;
        ChannelMessage t;
        t <- mod_1783.get(0);
        mod_1784.put(0, t);
    endrule
    rule rule_2321;
        ChannelMessage t;
        t <- mod_1784.get(0);
        mod_1783.put(1, t);
    endrule
    rule rule_2322;
        ChannelMessage t;
        t <- mod_1790.get(0);
        mod_1789.put(0, t);
    endrule
    rule rule_2323;
        ChannelMessage t;
        t <- mod_1779.get(0);
        mod_1781.put(0, t);
    endrule
    rule rule_2324;
        ChannelMessage t;
        t <- mod_1770.get(0);
        mod_1795.put(0, t);
    endrule
    rule rule_2325;
        ChannelMessage t;
        t <- mod_1770.get(1);
        mod_1771.put(0, t);
    endrule
    rule rule_2326;
        ChannelMessage t;
        t <- mod_1775.get(1);
        mod_1776.put(0, t);
    endrule
    rule rule_2327;
        ChannelMessage t;
        t <- mod_1785.get(0);
        mod_1783.put(0, t);
    endrule
    rule rule_2328;
        ChannelMessage t;
        t <- mod_1802.get(0);
        mod_1769.put(1, t);
    endrule
    rule rule_2329;
        ChannelMessage t;
        t <- mod_1803.get(1);
        mod_1767.put(1, t);
    endrule
    rule rule_2330;
        ChannelMessage t;
        t <- mod_1766.get(0);
        mod_1767.put(0, t);
    endrule
    rule rule_2331;
        ChannelMessage t;
        t <- mod_1778.get(0);
        mod_1782.put(0, t);
    endrule
    rule rule_2332;
        ChannelMessage t;
        t <- mod_1782.get(1);
        mod_1778.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1764.put(0, t);
        end
        if (i == 1) begin
            mod_1780.put(0, t);
        end
        if (i == 2) begin
            mod_1786.put(0, t);
        end
        if (i == 3) begin
            mod_1794.put(0, t);
        end
        if (i == 4) begin
            mod_1800.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_1768.get(0);
        end
        if (i == 2) begin
            t <- mod_1768.get(1);
        end
        if (i == 0) begin
            t <- mod_1768.get(2);
        end
        if (i == 1) begin
            t <- mod_1780.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6078 (Operation_IFC);
    Operation_IFC mod_1805_inner <- mkReshape(2, 64);
    Operation_IFC mod_1805 <- mkDebugOperation(mod_1805_inner, "mod_1805");
    Operation_IFC mod_1806_inner <- mkFlatten(1);
    Operation_IFC mod_1806 <- mkDebugOperation(mod_1806_inner, "mod_1806");
    Operation_IFC mod_1807_inner <- mkFlatten(2);
    Operation_IFC mod_1807 <- mkDebugOperation(mod_1807_inner, "mod_1807");
    Operation_IFC mod_1808_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1808 <- mkDebugOperation(mod_1808_inner, "mod_1808");
    Broadcast_IFC#(4) mod_1809_inner <- mkBroadcast(4);
    Operation_IFC mod_1809 <- mkDebugOperation(mod_1809_inner.op, "mod_1809");
    PMU_IFC mod_1810_bufferize <- mkPMU(2);
    Operation_IFC mod_1810_inner = mod_1810_bufferize.operation;
    Operation_IFC mod_1810 <- mkDebugOperation(mod_1810_inner, "mod_1810");
    Broadcast_IFC#(2) mod_1811_inner <- mkBroadcast(2);
    Operation_IFC mod_1811 <- mkDebugOperation(mod_1811_inner.op, "mod_1811");
    PMU_IFC mod_1812_bufferize <- mkPMU(1);
    Operation_IFC mod_1812_inner = mod_1812_bufferize.operation;
    Operation_IFC mod_1812 <- mkDebugOperation(mod_1812_inner, "mod_1812");
    Operation_IFC mod_1813_inner <- mkBinaryMap(1112, matmul_t_tile);
    Operation_IFC mod_1813 <- mkDebugOperation(mod_1813_inner, "mod_1813");
    Operation_IFC mod_1814_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1814 <- mkDebugOperation(mod_1814_inner, "mod_1814");
    Operation_IFC mod_1815_inner <- mkBinaryMap(1880, mul_tile);
    Operation_IFC mod_1815 <- mkDebugOperation(mod_1815_inner, "mod_1815");
    PMU_IFC mod_1816_bufferize <- mkPMU(1);
    Operation_IFC mod_1816_inner = mod_1816_bufferize.operation;
    Operation_IFC mod_1816 <- mkDebugOperation(mod_1816_inner, "mod_1816");
    Operation_IFC mod_1817_inner <- mkBinaryMap(2475, matmul_t_tile);
    Operation_IFC mod_1817 <- mkDebugOperation(mod_1817_inner, "mod_1817");
    Operation_IFC mod_1818_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1818 <- mkDebugOperation(mod_1818_inner, "mod_1818");
    Operation_IFC mod_1819_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1819 <- mkDebugOperation(mod_1819_inner, "mod_1819");
    Operation_IFC mod_1820_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1820 <- mkDebugOperation(mod_1820_inner, "mod_1820");
    Operation_IFC mod_1821_inner <- mkBinaryMap(2779, mul_tile);
    Operation_IFC mod_1821 <- mkDebugOperation(mod_1821_inner, "mod_1821");
    PMU_IFC mod_1822_bufferize <- mkPMU(1);
    Operation_IFC mod_1822_inner = mod_1822_bufferize.operation;
    Operation_IFC mod_1822 <- mkDebugOperation(mod_1822_inner, "mod_1822");
    PMU_IFC mod_1823_bufferize <- mkPMU(2);
    Operation_IFC mod_1823_inner = mod_1823_bufferize.operation;
    Operation_IFC mod_1823 <- mkDebugOperation(mod_1823_inner, "mod_1823");
    PMU_IFC mod_1824_bufferize <- mkPMU(2);
    Operation_IFC mod_1824_inner = mod_1824_bufferize.operation;
    Operation_IFC mod_1824 <- mkDebugOperation(mod_1824_inner, "mod_1824");
    Operation_IFC mod_1825_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1825 <- mkDebugOperation(mod_1825_inner, "mod_1825");
    Operation_IFC mod_1826_inner <- mkFlatten(1);
    Operation_IFC mod_1826 <- mkDebugOperation(mod_1826_inner, "mod_1826");
    Operation_IFC mod_1827_inner <- mkFlatten(0);
    Operation_IFC mod_1827 <- mkDebugOperation(mod_1827_inner, "mod_1827");
    Operation_IFC mod_1828_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1828 <- mkDebugOperation(mod_1828_inner, "mod_1828");
    Operation_IFC mod_1829_inner <- mkUnaryMap(1752, silu_tile);
    Operation_IFC mod_1829 <- mkDebugOperation(mod_1829_inner, "mod_1829");
    Operation_IFC mod_1830_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1830 <- mkDebugOperation(mod_1830_inner, "mod_1830");
    Operation_IFC mod_1831_inner <- mkBinaryMap(1624, matmul_t_tile);
    Operation_IFC mod_1831 <- mkDebugOperation(mod_1831_inner, "mod_1831");
    PMU_IFC mod_1832_bufferize <- mkPMU(2);
    Operation_IFC mod_1832_inner = mod_1832_bufferize.operation;
    Operation_IFC mod_1832 <- mkDebugOperation(mod_1832_inner, "mod_1832");
    Operation_IFC mod_1833_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1833 <- mkDebugOperation(mod_1833_inner, "mod_1833");
    Operation_IFC mod_1834_inner <- mkFlatten(1);
    Operation_IFC mod_1834 <- mkDebugOperation(mod_1834_inner, "mod_1834");
    Operation_IFC mod_1835_inner <- mkFlatten(0);
    Operation_IFC mod_1835 <- mkDebugOperation(mod_1835_inner, "mod_1835");
    PMU_IFC mod_1836_bufferize <- mkPMU(1);
    Operation_IFC mod_1836_inner = mod_1836_bufferize.operation;
    Operation_IFC mod_1836 <- mkDebugOperation(mod_1836_inner, "mod_1836");
    Operation_IFC mod_1837_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1837 <- mkDebugOperation(mod_1837_inner, "mod_1837");
    PMU_IFC mod_1838_bufferize <- mkPMU(2);
    Operation_IFC mod_1838_inner = mod_1838_bufferize.operation;
    Operation_IFC mod_1838 <- mkDebugOperation(mod_1838_inner, "mod_1838");
    Operation_IFC mod_1839_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1839 <- mkDebugOperation(mod_1839_inner, "mod_1839");
    Operation_IFC mod_1840_inner <- mkFlatten(1);
    Operation_IFC mod_1840 <- mkDebugOperation(mod_1840_inner, "mod_1840");
    Operation_IFC mod_1841_inner <- mkFlatten(0);
    Operation_IFC mod_1841 <- mkDebugOperation(mod_1841_inner, "mod_1841");
    Operation_IFC mod_1842_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1842 <- mkDebugOperation(mod_1842_inner, "mod_1842");
    Operation_IFC mod_1843_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1843 <- mkDebugOperation(mod_1843_inner, "mod_1843");
    PMU_IFC mod_1844_bufferize <- mkPMU(2);
    Operation_IFC mod_1844_inner = mod_1844_bufferize.operation;
    Operation_IFC mod_1844 <- mkDebugOperation(mod_1844_inner, "mod_1844");
    rule rule_2333;
        ChannelMessage t;
        t <- mod_1813.get(0);
        mod_1814.put(0, t);
    endrule
    rule rule_2334;
        ChannelMessage t;
        t <- mod_1828.get(0);
        mod_1816.put(1, t);
    endrule
    rule rule_2335;
        ChannelMessage t;
        t <- mod_1808.get(0);
        mod_1844.put(0, t);
    endrule
    rule rule_2336;
        ChannelMessage t;
        t <- mod_1834.get(0);
        mod_1832.put(0, t);
    endrule
    rule rule_2337;
        ChannelMessage t;
        t <- mod_1839.get(0);
        mod_1838.put(1, t);
    endrule
    rule rule_2338;
        ChannelMessage t;
        t <- mod_1805.get(0);
        mod_1806.put(0, t);
    endrule
    rule rule_2339;
        ChannelMessage t;
        t <- mod_1826.get(0);
        mod_1824.put(0, t);
    endrule
    rule rule_2340;
        ChannelMessage t;
        t <- mod_1808.get(1);
        mod_1809.put(0, t);
    endrule
    rule rule_2341;
        ChannelMessage t;
        t <- mod_1824.get(1);
        mod_1817.put(1, t);
    endrule
    rule rule_2342;
        ChannelMessage t;
        t <- mod_1822.get(1);
        mod_1820.put(1, t);
    endrule
    rule rule_2343;
        ChannelMessage t;
        t <- mod_1815.get(0);
        mod_1816.put(0, t);
    endrule
    rule rule_2344;
        ChannelMessage t;
        t <- mod_1812.get(1);
        mod_1813.put(0, t);
    endrule
    rule rule_2345;
        ChannelMessage t;
        t <- mod_1818.get(0);
        mod_1819.put(0, t);
    endrule
    rule rule_2346;
        ChannelMessage t;
        t <- mod_1831.get(0);
        mod_1830.put(0, t);
    endrule
    rule rule_2347;
        ChannelMessage t;
        t <- mod_1806.get(0);
        mod_1807.put(0, t);
    endrule
    rule rule_2348;
        ChannelMessage t;
        t <- mod_1835.get(0);
        mod_1834.put(0, t);
    endrule
    rule rule_2349;
        ChannelMessage t;
        t <- mod_1823.get(0);
        mod_1823.put(1, t);
    endrule
    rule rule_2350;
        ChannelMessage t;
        t <- mod_1832.get(0);
        mod_1833.put(0, t);
    endrule
    rule rule_2351;
        ChannelMessage t;
        t <- mod_1812.get(0);
        mod_1842.put(0, t);
    endrule
    rule rule_2352;
        ChannelMessage t;
        t <- mod_1838.get(0);
        mod_1839.put(0, t);
    endrule
    rule rule_2353;
        ChannelMessage t;
        t <- mod_1811.get(0);
        mod_1836.put(0, t);
    endrule
    rule rule_2354;
        ChannelMessage t;
        t <- mod_1838.get(1);
        mod_1813.put(1, t);
    endrule
    rule rule_2355;
        ChannelMessage t;
        t <- mod_1832.get(1);
        mod_1831.put(1, t);
    endrule
    rule rule_2356;
        ChannelMessage t;
        t <- mod_1809.get(3);
        mod_1810.put(0, t);
    endrule
    rule rule_2357;
        ChannelMessage t;
        t <- mod_1816.get(0);
        mod_1828.put(0, t);
    endrule
    rule rule_2358;
        ChannelMessage t;
        t <- mod_1827.get(0);
        mod_1826.put(0, t);
    endrule
    rule rule_2359;
        ChannelMessage t;
        t <- mod_1810.get(0);
        mod_1843.put(0, t);
    endrule
    rule rule_2360;
        ChannelMessage t;
        t <- mod_1823.get(1);
        mod_1819.put(1, t);
    endrule
    rule rule_2361;
        ChannelMessage t;
        t <- mod_1836.get(0);
        mod_1837.put(0, t);
    endrule
    rule rule_2362;
        ChannelMessage t;
        t <- mod_1811.get(1);
        mod_1812.put(0, t);
    endrule
    rule rule_2363;
        ChannelMessage t;
        t <- mod_1814.get(0);
        mod_1815.put(0, t);
    endrule
    rule rule_2364;
        ChannelMessage t;
        t <- mod_1825.get(0);
        mod_1824.put(1, t);
    endrule
    rule rule_2365;
        ChannelMessage t;
        t <- mod_1824.get(0);
        mod_1825.put(0, t);
    endrule
    rule rule_2366;
        ChannelMessage t;
        t <- mod_1817.get(0);
        mod_1818.put(0, t);
    endrule
    rule rule_2367;
        ChannelMessage t;
        t <- mod_1819.get(0);
        mod_1823.put(0, t);
    endrule
    rule rule_2368;
        ChannelMessage t;
        t <- mod_1820.get(0);
        mod_1822.put(0, t);
    endrule
    rule rule_2369;
        ChannelMessage t;
        t <- mod_1819.get(1);
        mod_1820.put(0, t);
    endrule
    rule rule_2370;
        ChannelMessage t;
        t <- mod_1807.get(0);
        mod_1808.put(0, t);
    endrule
    rule rule_2371;
        ChannelMessage t;
        t <- mod_1829.get(0);
        mod_1815.put(1, t);
    endrule
    rule rule_2372;
        ChannelMessage t;
        t <- mod_1836.get(1);
        mod_1831.put(0, t);
    endrule
    rule rule_2373;
        ChannelMessage t;
        t <- mod_1842.get(0);
        mod_1812.put(1, t);
    endrule
    rule rule_2374;
        ChannelMessage t;
        t <- mod_1810.get(1);
        mod_1811.put(0, t);
    endrule
    rule rule_2375;
        ChannelMessage t;
        t <- mod_1837.get(0);
        mod_1836.put(1, t);
    endrule
    rule rule_2376;
        ChannelMessage t;
        t <- mod_1816.get(1);
        mod_1817.put(0, t);
    endrule
    rule rule_2377;
        ChannelMessage t;
        t <- mod_1822.get(0);
        mod_1822.put(1, t);
    endrule
    rule rule_2378;
        ChannelMessage t;
        t <- mod_1833.get(0);
        mod_1832.put(1, t);
    endrule
    rule rule_2379;
        ChannelMessage t;
        t <- mod_1820.get(1);
        mod_1821.put(1, t);
    endrule
    rule rule_2380;
        ChannelMessage t;
        t <- mod_1841.get(0);
        mod_1840.put(0, t);
    endrule
    rule rule_2381;
        ChannelMessage t;
        t <- mod_1843.get(0);
        mod_1810.put(1, t);
    endrule
    rule rule_2382;
        ChannelMessage t;
        t <- mod_1844.get(0);
        mod_1844.put(1, t);
    endrule
    rule rule_2383;
        ChannelMessage t;
        t <- mod_1844.get(1);
        mod_1808.put(1, t);
    endrule
    rule rule_2384;
        ChannelMessage t;
        t <- mod_1840.get(0);
        mod_1838.put(0, t);
    endrule
    rule rule_2385;
        ChannelMessage t;
        t <- mod_1830.get(0);
        mod_1829.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1805.put(0, t);
        end
        if (i == 1) begin
            mod_1821.put(0, t);
        end
        if (i == 2) begin
            mod_1827.put(0, t);
        end
        if (i == 3) begin
            mod_1835.put(0, t);
        end
        if (i == 4) begin
            mod_1841.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_1809.get(0);
        end
        if (i == 1) begin
            t <- mod_1809.get(1);
        end
        if (i == 0) begin
            t <- mod_1809.get(2);
        end
        if (i == 2) begin
            t <- mod_1821.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6079 (Operation_IFC);
    Operation_IFC mod_1846_inner <- mkReshape(2, 64);
    Operation_IFC mod_1846 <- mkDebugOperation(mod_1846_inner, "mod_1846");
    Operation_IFC mod_1847_inner <- mkFlatten(1);
    Operation_IFC mod_1847 <- mkDebugOperation(mod_1847_inner, "mod_1847");
    Operation_IFC mod_1848_inner <- mkFlatten(2);
    Operation_IFC mod_1848 <- mkDebugOperation(mod_1848_inner, "mod_1848");
    Operation_IFC mod_1849_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1849 <- mkDebugOperation(mod_1849_inner, "mod_1849");
    Broadcast_IFC#(4) mod_1850_inner <- mkBroadcast(4);
    Operation_IFC mod_1850 <- mkDebugOperation(mod_1850_inner.op, "mod_1850");
    PMU_IFC mod_1851_bufferize <- mkPMU(2);
    Operation_IFC mod_1851_inner = mod_1851_bufferize.operation;
    Operation_IFC mod_1851 <- mkDebugOperation(mod_1851_inner, "mod_1851");
    Broadcast_IFC#(2) mod_1852_inner <- mkBroadcast(2);
    Operation_IFC mod_1852 <- mkDebugOperation(mod_1852_inner.op, "mod_1852");
    PMU_IFC mod_1853_bufferize <- mkPMU(1);
    Operation_IFC mod_1853_inner = mod_1853_bufferize.operation;
    Operation_IFC mod_1853 <- mkDebugOperation(mod_1853_inner, "mod_1853");
    Operation_IFC mod_1854_inner <- mkBinaryMap(1111, matmul_t_tile);
    Operation_IFC mod_1854 <- mkDebugOperation(mod_1854_inner, "mod_1854");
    Operation_IFC mod_1855_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1855 <- mkDebugOperation(mod_1855_inner, "mod_1855");
    Operation_IFC mod_1856_inner <- mkBinaryMap(1879, mul_tile);
    Operation_IFC mod_1856 <- mkDebugOperation(mod_1856_inner, "mod_1856");
    PMU_IFC mod_1857_bufferize <- mkPMU(1);
    Operation_IFC mod_1857_inner = mod_1857_bufferize.operation;
    Operation_IFC mod_1857 <- mkDebugOperation(mod_1857_inner, "mod_1857");
    Operation_IFC mod_1858_inner <- mkBinaryMap(2473, matmul_t_tile);
    Operation_IFC mod_1858 <- mkDebugOperation(mod_1858_inner, "mod_1858");
    Operation_IFC mod_1859_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1859 <- mkDebugOperation(mod_1859_inner, "mod_1859");
    Operation_IFC mod_1860_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1860 <- mkDebugOperation(mod_1860_inner, "mod_1860");
    Operation_IFC mod_1861_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1861 <- mkDebugOperation(mod_1861_inner, "mod_1861");
    Operation_IFC mod_1862_inner <- mkBinaryMap(2778, mul_tile);
    Operation_IFC mod_1862 <- mkDebugOperation(mod_1862_inner, "mod_1862");
    PMU_IFC mod_1863_bufferize <- mkPMU(1);
    Operation_IFC mod_1863_inner = mod_1863_bufferize.operation;
    Operation_IFC mod_1863 <- mkDebugOperation(mod_1863_inner, "mod_1863");
    PMU_IFC mod_1864_bufferize <- mkPMU(2);
    Operation_IFC mod_1864_inner = mod_1864_bufferize.operation;
    Operation_IFC mod_1864 <- mkDebugOperation(mod_1864_inner, "mod_1864");
    PMU_IFC mod_1865_bufferize <- mkPMU(2);
    Operation_IFC mod_1865_inner = mod_1865_bufferize.operation;
    Operation_IFC mod_1865 <- mkDebugOperation(mod_1865_inner, "mod_1865");
    Operation_IFC mod_1866_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1866 <- mkDebugOperation(mod_1866_inner, "mod_1866");
    Operation_IFC mod_1867_inner <- mkFlatten(1);
    Operation_IFC mod_1867 <- mkDebugOperation(mod_1867_inner, "mod_1867");
    Operation_IFC mod_1868_inner <- mkFlatten(0);
    Operation_IFC mod_1868 <- mkDebugOperation(mod_1868_inner, "mod_1868");
    Operation_IFC mod_1869_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1869 <- mkDebugOperation(mod_1869_inner, "mod_1869");
    Operation_IFC mod_1870_inner <- mkUnaryMap(1751, silu_tile);
    Operation_IFC mod_1870 <- mkDebugOperation(mod_1870_inner, "mod_1870");
    Operation_IFC mod_1871_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1871 <- mkDebugOperation(mod_1871_inner, "mod_1871");
    Operation_IFC mod_1872_inner <- mkBinaryMap(1623, matmul_t_tile);
    Operation_IFC mod_1872 <- mkDebugOperation(mod_1872_inner, "mod_1872");
    PMU_IFC mod_1873_bufferize <- mkPMU(2);
    Operation_IFC mod_1873_inner = mod_1873_bufferize.operation;
    Operation_IFC mod_1873 <- mkDebugOperation(mod_1873_inner, "mod_1873");
    Operation_IFC mod_1874_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1874 <- mkDebugOperation(mod_1874_inner, "mod_1874");
    Operation_IFC mod_1875_inner <- mkFlatten(1);
    Operation_IFC mod_1875 <- mkDebugOperation(mod_1875_inner, "mod_1875");
    Operation_IFC mod_1876_inner <- mkFlatten(0);
    Operation_IFC mod_1876 <- mkDebugOperation(mod_1876_inner, "mod_1876");
    PMU_IFC mod_1877_bufferize <- mkPMU(1);
    Operation_IFC mod_1877_inner = mod_1877_bufferize.operation;
    Operation_IFC mod_1877 <- mkDebugOperation(mod_1877_inner, "mod_1877");
    Operation_IFC mod_1878_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1878 <- mkDebugOperation(mod_1878_inner, "mod_1878");
    PMU_IFC mod_1879_bufferize <- mkPMU(2);
    Operation_IFC mod_1879_inner = mod_1879_bufferize.operation;
    Operation_IFC mod_1879 <- mkDebugOperation(mod_1879_inner, "mod_1879");
    Operation_IFC mod_1880_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1880 <- mkDebugOperation(mod_1880_inner, "mod_1880");
    Operation_IFC mod_1881_inner <- mkFlatten(1);
    Operation_IFC mod_1881 <- mkDebugOperation(mod_1881_inner, "mod_1881");
    Operation_IFC mod_1882_inner <- mkFlatten(0);
    Operation_IFC mod_1882 <- mkDebugOperation(mod_1882_inner, "mod_1882");
    Operation_IFC mod_1883_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1883 <- mkDebugOperation(mod_1883_inner, "mod_1883");
    Operation_IFC mod_1884_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1884 <- mkDebugOperation(mod_1884_inner, "mod_1884");
    PMU_IFC mod_1885_bufferize <- mkPMU(2);
    Operation_IFC mod_1885_inner = mod_1885_bufferize.operation;
    Operation_IFC mod_1885 <- mkDebugOperation(mod_1885_inner, "mod_1885");
    rule rule_2386;
        ChannelMessage t;
        t <- mod_1859.get(0);
        mod_1860.put(0, t);
    endrule
    rule rule_2387;
        ChannelMessage t;
        t <- mod_1855.get(0);
        mod_1856.put(0, t);
    endrule
    rule rule_2388;
        ChannelMessage t;
        t <- mod_1860.get(1);
        mod_1861.put(0, t);
    endrule
    rule rule_2389;
        ChannelMessage t;
        t <- mod_1863.get(0);
        mod_1863.put(1, t);
    endrule
    rule rule_2390;
        ChannelMessage t;
        t <- mod_1873.get(1);
        mod_1872.put(1, t);
    endrule
    rule rule_2391;
        ChannelMessage t;
        t <- mod_1864.get(0);
        mod_1864.put(1, t);
    endrule
    rule rule_2392;
        ChannelMessage t;
        t <- mod_1851.get(0);
        mod_1884.put(0, t);
    endrule
    rule rule_2393;
        ChannelMessage t;
        t <- mod_1877.get(1);
        mod_1872.put(0, t);
    endrule
    rule rule_2394;
        ChannelMessage t;
        t <- mod_1871.get(0);
        mod_1870.put(0, t);
    endrule
    rule rule_2395;
        ChannelMessage t;
        t <- mod_1868.get(0);
        mod_1867.put(0, t);
    endrule
    rule rule_2396;
        ChannelMessage t;
        t <- mod_1864.get(1);
        mod_1860.put(1, t);
    endrule
    rule rule_2397;
        ChannelMessage t;
        t <- mod_1870.get(0);
        mod_1856.put(1, t);
    endrule
    rule rule_2398;
        ChannelMessage t;
        t <- mod_1866.get(0);
        mod_1865.put(1, t);
    endrule
    rule rule_2399;
        ChannelMessage t;
        t <- mod_1861.get(1);
        mod_1862.put(1, t);
    endrule
    rule rule_2400;
        ChannelMessage t;
        t <- mod_1856.get(0);
        mod_1857.put(0, t);
    endrule
    rule rule_2401;
        ChannelMessage t;
        t <- mod_1865.get(1);
        mod_1858.put(1, t);
    endrule
    rule rule_2402;
        ChannelMessage t;
        t <- mod_1857.get(0);
        mod_1869.put(0, t);
    endrule
    rule rule_2403;
        ChannelMessage t;
        t <- mod_1854.get(0);
        mod_1855.put(0, t);
    endrule
    rule rule_2404;
        ChannelMessage t;
        t <- mod_1857.get(1);
        mod_1858.put(0, t);
    endrule
    rule rule_2405;
        ChannelMessage t;
        t <- mod_1881.get(0);
        mod_1879.put(0, t);
    endrule
    rule rule_2406;
        ChannelMessage t;
        t <- mod_1878.get(0);
        mod_1877.put(1, t);
    endrule
    rule rule_2407;
        ChannelMessage t;
        t <- mod_1876.get(0);
        mod_1875.put(0, t);
    endrule
    rule rule_2408;
        ChannelMessage t;
        t <- mod_1852.get(0);
        mod_1877.put(0, t);
    endrule
    rule rule_2409;
        ChannelMessage t;
        t <- mod_1851.get(1);
        mod_1852.put(0, t);
    endrule
    rule rule_2410;
        ChannelMessage t;
        t <- mod_1863.get(1);
        mod_1861.put(1, t);
    endrule
    rule rule_2411;
        ChannelMessage t;
        t <- mod_1869.get(0);
        mod_1857.put(1, t);
    endrule
    rule rule_2412;
        ChannelMessage t;
        t <- mod_1867.get(0);
        mod_1865.put(0, t);
    endrule
    rule rule_2413;
        ChannelMessage t;
        t <- mod_1847.get(0);
        mod_1848.put(0, t);
    endrule
    rule rule_2414;
        ChannelMessage t;
        t <- mod_1849.get(0);
        mod_1885.put(0, t);
    endrule
    rule rule_2415;
        ChannelMessage t;
        t <- mod_1865.get(0);
        mod_1866.put(0, t);
    endrule
    rule rule_2416;
        ChannelMessage t;
        t <- mod_1875.get(0);
        mod_1873.put(0, t);
    endrule
    rule rule_2417;
        ChannelMessage t;
        t <- mod_1850.get(3);
        mod_1851.put(0, t);
    endrule
    rule rule_2418;
        ChannelMessage t;
        t <- mod_1848.get(0);
        mod_1849.put(0, t);
    endrule
    rule rule_2419;
        ChannelMessage t;
        t <- mod_1872.get(0);
        mod_1871.put(0, t);
    endrule
    rule rule_2420;
        ChannelMessage t;
        t <- mod_1882.get(0);
        mod_1881.put(0, t);
    endrule
    rule rule_2421;
        ChannelMessage t;
        t <- mod_1853.get(1);
        mod_1854.put(0, t);
    endrule
    rule rule_2422;
        ChannelMessage t;
        t <- mod_1883.get(0);
        mod_1853.put(1, t);
    endrule
    rule rule_2423;
        ChannelMessage t;
        t <- mod_1885.get(0);
        mod_1885.put(1, t);
    endrule
    rule rule_2424;
        ChannelMessage t;
        t <- mod_1849.get(1);
        mod_1850.put(0, t);
    endrule
    rule rule_2425;
        ChannelMessage t;
        t <- mod_1879.get(1);
        mod_1854.put(1, t);
    endrule
    rule rule_2426;
        ChannelMessage t;
        t <- mod_1877.get(0);
        mod_1878.put(0, t);
    endrule
    rule rule_2427;
        ChannelMessage t;
        t <- mod_1873.get(0);
        mod_1874.put(0, t);
    endrule
    rule rule_2428;
        ChannelMessage t;
        t <- mod_1874.get(0);
        mod_1873.put(1, t);
    endrule
    rule rule_2429;
        ChannelMessage t;
        t <- mod_1852.get(1);
        mod_1853.put(0, t);
    endrule
    rule rule_2430;
        ChannelMessage t;
        t <- mod_1879.get(0);
        mod_1880.put(0, t);
    endrule
    rule rule_2431;
        ChannelMessage t;
        t <- mod_1860.get(0);
        mod_1864.put(0, t);
    endrule
    rule rule_2432;
        ChannelMessage t;
        t <- mod_1880.get(0);
        mod_1879.put(1, t);
    endrule
    rule rule_2433;
        ChannelMessage t;
        t <- mod_1861.get(0);
        mod_1863.put(0, t);
    endrule
    rule rule_2434;
        ChannelMessage t;
        t <- mod_1858.get(0);
        mod_1859.put(0, t);
    endrule
    rule rule_2435;
        ChannelMessage t;
        t <- mod_1846.get(0);
        mod_1847.put(0, t);
    endrule
    rule rule_2436;
        ChannelMessage t;
        t <- mod_1853.get(0);
        mod_1883.put(0, t);
    endrule
    rule rule_2437;
        ChannelMessage t;
        t <- mod_1884.get(0);
        mod_1851.put(1, t);
    endrule
    rule rule_2438;
        ChannelMessage t;
        t <- mod_1885.get(1);
        mod_1849.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1846.put(0, t);
        end
        if (i == 1) begin
            mod_1862.put(0, t);
        end
        if (i == 2) begin
            mod_1868.put(0, t);
        end
        if (i == 3) begin
            mod_1876.put(0, t);
        end
        if (i == 4) begin
            mod_1882.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_1850.get(0);
        end
        if (i == 2) begin
            t <- mod_1850.get(1);
        end
        if (i == 3) begin
            t <- mod_1850.get(2);
        end
        if (i == 0) begin
            t <- mod_1862.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6080 (Operation_IFC);
    Operation_IFC mod_1887_inner <- mkReshape(2, 64);
    Operation_IFC mod_1887 <- mkDebugOperation(mod_1887_inner, "mod_1887");
    Operation_IFC mod_1888_inner <- mkFlatten(1);
    Operation_IFC mod_1888 <- mkDebugOperation(mod_1888_inner, "mod_1888");
    Operation_IFC mod_1889_inner <- mkFlatten(2);
    Operation_IFC mod_1889 <- mkDebugOperation(mod_1889_inner, "mod_1889");
    Operation_IFC mod_1890_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1890 <- mkDebugOperation(mod_1890_inner, "mod_1890");
    Broadcast_IFC#(4) mod_1891_inner <- mkBroadcast(4);
    Operation_IFC mod_1891 <- mkDebugOperation(mod_1891_inner.op, "mod_1891");
    PMU_IFC mod_1892_bufferize <- mkPMU(2);
    Operation_IFC mod_1892_inner = mod_1892_bufferize.operation;
    Operation_IFC mod_1892 <- mkDebugOperation(mod_1892_inner, "mod_1892");
    Broadcast_IFC#(2) mod_1893_inner <- mkBroadcast(2);
    Operation_IFC mod_1893 <- mkDebugOperation(mod_1893_inner.op, "mod_1893");
    PMU_IFC mod_1894_bufferize <- mkPMU(1);
    Operation_IFC mod_1894_inner = mod_1894_bufferize.operation;
    Operation_IFC mod_1894 <- mkDebugOperation(mod_1894_inner, "mod_1894");
    Operation_IFC mod_1895_inner <- mkBinaryMap(1110, matmul_t_tile);
    Operation_IFC mod_1895 <- mkDebugOperation(mod_1895_inner, "mod_1895");
    Operation_IFC mod_1896_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1896 <- mkDebugOperation(mod_1896_inner, "mod_1896");
    Operation_IFC mod_1897_inner <- mkBinaryMap(1878, mul_tile);
    Operation_IFC mod_1897 <- mkDebugOperation(mod_1897_inner, "mod_1897");
    PMU_IFC mod_1898_bufferize <- mkPMU(1);
    Operation_IFC mod_1898_inner = mod_1898_bufferize.operation;
    Operation_IFC mod_1898 <- mkDebugOperation(mod_1898_inner, "mod_1898");
    Operation_IFC mod_1899_inner <- mkBinaryMap(2471, matmul_t_tile);
    Operation_IFC mod_1899 <- mkDebugOperation(mod_1899_inner, "mod_1899");
    Operation_IFC mod_1900_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1900 <- mkDebugOperation(mod_1900_inner, "mod_1900");
    Operation_IFC mod_1901_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1901 <- mkDebugOperation(mod_1901_inner, "mod_1901");
    Operation_IFC mod_1902_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1902 <- mkDebugOperation(mod_1902_inner, "mod_1902");
    Operation_IFC mod_1903_inner <- mkBinaryMap(2777, mul_tile);
    Operation_IFC mod_1903 <- mkDebugOperation(mod_1903_inner, "mod_1903");
    PMU_IFC mod_1904_bufferize <- mkPMU(1);
    Operation_IFC mod_1904_inner = mod_1904_bufferize.operation;
    Operation_IFC mod_1904 <- mkDebugOperation(mod_1904_inner, "mod_1904");
    PMU_IFC mod_1905_bufferize <- mkPMU(2);
    Operation_IFC mod_1905_inner = mod_1905_bufferize.operation;
    Operation_IFC mod_1905 <- mkDebugOperation(mod_1905_inner, "mod_1905");
    PMU_IFC mod_1906_bufferize <- mkPMU(2);
    Operation_IFC mod_1906_inner = mod_1906_bufferize.operation;
    Operation_IFC mod_1906 <- mkDebugOperation(mod_1906_inner, "mod_1906");
    Operation_IFC mod_1907_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1907 <- mkDebugOperation(mod_1907_inner, "mod_1907");
    Operation_IFC mod_1908_inner <- mkFlatten(1);
    Operation_IFC mod_1908 <- mkDebugOperation(mod_1908_inner, "mod_1908");
    Operation_IFC mod_1909_inner <- mkFlatten(0);
    Operation_IFC mod_1909 <- mkDebugOperation(mod_1909_inner, "mod_1909");
    Operation_IFC mod_1910_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1910 <- mkDebugOperation(mod_1910_inner, "mod_1910");
    Operation_IFC mod_1911_inner <- mkUnaryMap(1750, silu_tile);
    Operation_IFC mod_1911 <- mkDebugOperation(mod_1911_inner, "mod_1911");
    Operation_IFC mod_1912_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1912 <- mkDebugOperation(mod_1912_inner, "mod_1912");
    Operation_IFC mod_1913_inner <- mkBinaryMap(1622, matmul_t_tile);
    Operation_IFC mod_1913 <- mkDebugOperation(mod_1913_inner, "mod_1913");
    PMU_IFC mod_1914_bufferize <- mkPMU(2);
    Operation_IFC mod_1914_inner = mod_1914_bufferize.operation;
    Operation_IFC mod_1914 <- mkDebugOperation(mod_1914_inner, "mod_1914");
    Operation_IFC mod_1915_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1915 <- mkDebugOperation(mod_1915_inner, "mod_1915");
    Operation_IFC mod_1916_inner <- mkFlatten(1);
    Operation_IFC mod_1916 <- mkDebugOperation(mod_1916_inner, "mod_1916");
    Operation_IFC mod_1917_inner <- mkFlatten(0);
    Operation_IFC mod_1917 <- mkDebugOperation(mod_1917_inner, "mod_1917");
    PMU_IFC mod_1918_bufferize <- mkPMU(1);
    Operation_IFC mod_1918_inner = mod_1918_bufferize.operation;
    Operation_IFC mod_1918 <- mkDebugOperation(mod_1918_inner, "mod_1918");
    Operation_IFC mod_1919_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1919 <- mkDebugOperation(mod_1919_inner, "mod_1919");
    PMU_IFC mod_1920_bufferize <- mkPMU(2);
    Operation_IFC mod_1920_inner = mod_1920_bufferize.operation;
    Operation_IFC mod_1920 <- mkDebugOperation(mod_1920_inner, "mod_1920");
    Operation_IFC mod_1921_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1921 <- mkDebugOperation(mod_1921_inner, "mod_1921");
    Operation_IFC mod_1922_inner <- mkFlatten(1);
    Operation_IFC mod_1922 <- mkDebugOperation(mod_1922_inner, "mod_1922");
    Operation_IFC mod_1923_inner <- mkFlatten(0);
    Operation_IFC mod_1923 <- mkDebugOperation(mod_1923_inner, "mod_1923");
    Operation_IFC mod_1924_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1924 <- mkDebugOperation(mod_1924_inner, "mod_1924");
    Operation_IFC mod_1925_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1925 <- mkDebugOperation(mod_1925_inner, "mod_1925");
    PMU_IFC mod_1926_bufferize <- mkPMU(2);
    Operation_IFC mod_1926_inner = mod_1926_bufferize.operation;
    Operation_IFC mod_1926 <- mkDebugOperation(mod_1926_inner, "mod_1926");
    rule rule_2439;
        ChannelMessage t;
        t <- mod_1926.get(0);
        mod_1926.put(1, t);
    endrule
    rule rule_2440;
        ChannelMessage t;
        t <- mod_1902.get(1);
        mod_1903.put(1, t);
    endrule
    rule rule_2441;
        ChannelMessage t;
        t <- mod_1891.get(3);
        mod_1892.put(0, t);
    endrule
    rule rule_2442;
        ChannelMessage t;
        t <- mod_1918.get(0);
        mod_1919.put(0, t);
    endrule
    rule rule_2443;
        ChannelMessage t;
        t <- mod_1904.get(0);
        mod_1904.put(1, t);
    endrule
    rule rule_2444;
        ChannelMessage t;
        t <- mod_1909.get(0);
        mod_1908.put(0, t);
    endrule
    rule rule_2445;
        ChannelMessage t;
        t <- mod_1896.get(0);
        mod_1897.put(0, t);
    endrule
    rule rule_2446;
        ChannelMessage t;
        t <- mod_1907.get(0);
        mod_1906.put(1, t);
    endrule
    rule rule_2447;
        ChannelMessage t;
        t <- mod_1914.get(1);
        mod_1913.put(1, t);
    endrule
    rule rule_2448;
        ChannelMessage t;
        t <- mod_1923.get(0);
        mod_1922.put(0, t);
    endrule
    rule rule_2449;
        ChannelMessage t;
        t <- mod_1887.get(0);
        mod_1888.put(0, t);
    endrule
    rule rule_2450;
        ChannelMessage t;
        t <- mod_1908.get(0);
        mod_1906.put(0, t);
    endrule
    rule rule_2451;
        ChannelMessage t;
        t <- mod_1914.get(0);
        mod_1915.put(0, t);
    endrule
    rule rule_2452;
        ChannelMessage t;
        t <- mod_1912.get(0);
        mod_1911.put(0, t);
    endrule
    rule rule_2453;
        ChannelMessage t;
        t <- mod_1899.get(0);
        mod_1900.put(0, t);
    endrule
    rule rule_2454;
        ChannelMessage t;
        t <- mod_1895.get(0);
        mod_1896.put(0, t);
    endrule
    rule rule_2455;
        ChannelMessage t;
        t <- mod_1898.get(1);
        mod_1899.put(0, t);
    endrule
    rule rule_2456;
        ChannelMessage t;
        t <- mod_1902.get(0);
        mod_1904.put(0, t);
    endrule
    rule rule_2457;
        ChannelMessage t;
        t <- mod_1925.get(0);
        mod_1892.put(1, t);
    endrule
    rule rule_2458;
        ChannelMessage t;
        t <- mod_1893.get(1);
        mod_1894.put(0, t);
    endrule
    rule rule_2459;
        ChannelMessage t;
        t <- mod_1922.get(0);
        mod_1920.put(0, t);
    endrule
    rule rule_2460;
        ChannelMessage t;
        t <- mod_1921.get(0);
        mod_1920.put(1, t);
    endrule
    rule rule_2461;
        ChannelMessage t;
        t <- mod_1889.get(0);
        mod_1890.put(0, t);
    endrule
    rule rule_2462;
        ChannelMessage t;
        t <- mod_1901.get(1);
        mod_1902.put(0, t);
    endrule
    rule rule_2463;
        ChannelMessage t;
        t <- mod_1920.get(1);
        mod_1895.put(1, t);
    endrule
    rule rule_2464;
        ChannelMessage t;
        t <- mod_1900.get(0);
        mod_1901.put(0, t);
    endrule
    rule rule_2465;
        ChannelMessage t;
        t <- mod_1897.get(0);
        mod_1898.put(0, t);
    endrule
    rule rule_2466;
        ChannelMessage t;
        t <- mod_1905.get(0);
        mod_1905.put(1, t);
    endrule
    rule rule_2467;
        ChannelMessage t;
        t <- mod_1892.get(0);
        mod_1925.put(0, t);
    endrule
    rule rule_2468;
        ChannelMessage t;
        t <- mod_1904.get(1);
        mod_1902.put(1, t);
    endrule
    rule rule_2469;
        ChannelMessage t;
        t <- mod_1926.get(1);
        mod_1890.put(1, t);
    endrule
    rule rule_2470;
        ChannelMessage t;
        t <- mod_1919.get(0);
        mod_1918.put(1, t);
    endrule
    rule rule_2471;
        ChannelMessage t;
        t <- mod_1920.get(0);
        mod_1921.put(0, t);
    endrule
    rule rule_2472;
        ChannelMessage t;
        t <- mod_1913.get(0);
        mod_1912.put(0, t);
    endrule
    rule rule_2473;
        ChannelMessage t;
        t <- mod_1905.get(1);
        mod_1901.put(1, t);
    endrule
    rule rule_2474;
        ChannelMessage t;
        t <- mod_1924.get(0);
        mod_1894.put(1, t);
    endrule
    rule rule_2475;
        ChannelMessage t;
        t <- mod_1890.get(0);
        mod_1926.put(0, t);
    endrule
    rule rule_2476;
        ChannelMessage t;
        t <- mod_1918.get(1);
        mod_1913.put(0, t);
    endrule
    rule rule_2477;
        ChannelMessage t;
        t <- mod_1901.get(0);
        mod_1905.put(0, t);
    endrule
    rule rule_2478;
        ChannelMessage t;
        t <- mod_1898.get(0);
        mod_1910.put(0, t);
    endrule
    rule rule_2479;
        ChannelMessage t;
        t <- mod_1906.get(0);
        mod_1907.put(0, t);
    endrule
    rule rule_2480;
        ChannelMessage t;
        t <- mod_1892.get(1);
        mod_1893.put(0, t);
    endrule
    rule rule_2481;
        ChannelMessage t;
        t <- mod_1915.get(0);
        mod_1914.put(1, t);
    endrule
    rule rule_2482;
        ChannelMessage t;
        t <- mod_1888.get(0);
        mod_1889.put(0, t);
    endrule
    rule rule_2483;
        ChannelMessage t;
        t <- mod_1917.get(0);
        mod_1916.put(0, t);
    endrule
    rule rule_2484;
        ChannelMessage t;
        t <- mod_1893.get(0);
        mod_1918.put(0, t);
    endrule
    rule rule_2485;
        ChannelMessage t;
        t <- mod_1906.get(1);
        mod_1899.put(1, t);
    endrule
    rule rule_2486;
        ChannelMessage t;
        t <- mod_1911.get(0);
        mod_1897.put(1, t);
    endrule
    rule rule_2487;
        ChannelMessage t;
        t <- mod_1894.get(1);
        mod_1895.put(0, t);
    endrule
    rule rule_2488;
        ChannelMessage t;
        t <- mod_1916.get(0);
        mod_1914.put(0, t);
    endrule
    rule rule_2489;
        ChannelMessage t;
        t <- mod_1894.get(0);
        mod_1924.put(0, t);
    endrule
    rule rule_2490;
        ChannelMessage t;
        t <- mod_1890.get(1);
        mod_1891.put(0, t);
    endrule
    rule rule_2491;
        ChannelMessage t;
        t <- mod_1910.get(0);
        mod_1898.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1887.put(0, t);
        end
        if (i == 1) begin
            mod_1903.put(0, t);
        end
        if (i == 2) begin
            mod_1909.put(0, t);
        end
        if (i == 3) begin
            mod_1917.put(0, t);
        end
        if (i == 4) begin
            mod_1923.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_1891.get(0);
        end
        if (i == 0) begin
            t <- mod_1891.get(1);
        end
        if (i == 3) begin
            t <- mod_1891.get(2);
        end
        if (i == 2) begin
            t <- mod_1903.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6081 (Operation_IFC);
    Operation_IFC mod_1928_inner <- mkReshape(2, 64);
    Operation_IFC mod_1928 <- mkDebugOperation(mod_1928_inner, "mod_1928");
    Operation_IFC mod_1929_inner <- mkFlatten(1);
    Operation_IFC mod_1929 <- mkDebugOperation(mod_1929_inner, "mod_1929");
    Operation_IFC mod_1930_inner <- mkFlatten(2);
    Operation_IFC mod_1930 <- mkDebugOperation(mod_1930_inner, "mod_1930");
    Operation_IFC mod_1931_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1931 <- mkDebugOperation(mod_1931_inner, "mod_1931");
    Broadcast_IFC#(4) mod_1932_inner <- mkBroadcast(4);
    Operation_IFC mod_1932 <- mkDebugOperation(mod_1932_inner.op, "mod_1932");
    PMU_IFC mod_1933_bufferize <- mkPMU(2);
    Operation_IFC mod_1933_inner = mod_1933_bufferize.operation;
    Operation_IFC mod_1933 <- mkDebugOperation(mod_1933_inner, "mod_1933");
    Broadcast_IFC#(2) mod_1934_inner <- mkBroadcast(2);
    Operation_IFC mod_1934 <- mkDebugOperation(mod_1934_inner.op, "mod_1934");
    PMU_IFC mod_1935_bufferize <- mkPMU(1);
    Operation_IFC mod_1935_inner = mod_1935_bufferize.operation;
    Operation_IFC mod_1935 <- mkDebugOperation(mod_1935_inner, "mod_1935");
    Operation_IFC mod_1936_inner <- mkBinaryMap(1109, matmul_t_tile);
    Operation_IFC mod_1936 <- mkDebugOperation(mod_1936_inner, "mod_1936");
    Operation_IFC mod_1937_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1937 <- mkDebugOperation(mod_1937_inner, "mod_1937");
    Operation_IFC mod_1938_inner <- mkBinaryMap(1877, mul_tile);
    Operation_IFC mod_1938 <- mkDebugOperation(mod_1938_inner, "mod_1938");
    PMU_IFC mod_1939_bufferize <- mkPMU(1);
    Operation_IFC mod_1939_inner = mod_1939_bufferize.operation;
    Operation_IFC mod_1939 <- mkDebugOperation(mod_1939_inner, "mod_1939");
    Operation_IFC mod_1940_inner <- mkBinaryMap(2469, matmul_t_tile);
    Operation_IFC mod_1940 <- mkDebugOperation(mod_1940_inner, "mod_1940");
    Operation_IFC mod_1941_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1941 <- mkDebugOperation(mod_1941_inner, "mod_1941");
    Operation_IFC mod_1942_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1942 <- mkDebugOperation(mod_1942_inner, "mod_1942");
    Operation_IFC mod_1943_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1943 <- mkDebugOperation(mod_1943_inner, "mod_1943");
    Operation_IFC mod_1944_inner <- mkBinaryMap(2776, mul_tile);
    Operation_IFC mod_1944 <- mkDebugOperation(mod_1944_inner, "mod_1944");
    PMU_IFC mod_1945_bufferize <- mkPMU(1);
    Operation_IFC mod_1945_inner = mod_1945_bufferize.operation;
    Operation_IFC mod_1945 <- mkDebugOperation(mod_1945_inner, "mod_1945");
    PMU_IFC mod_1946_bufferize <- mkPMU(2);
    Operation_IFC mod_1946_inner = mod_1946_bufferize.operation;
    Operation_IFC mod_1946 <- mkDebugOperation(mod_1946_inner, "mod_1946");
    PMU_IFC mod_1947_bufferize <- mkPMU(2);
    Operation_IFC mod_1947_inner = mod_1947_bufferize.operation;
    Operation_IFC mod_1947 <- mkDebugOperation(mod_1947_inner, "mod_1947");
    Operation_IFC mod_1948_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1948 <- mkDebugOperation(mod_1948_inner, "mod_1948");
    Operation_IFC mod_1949_inner <- mkFlatten(1);
    Operation_IFC mod_1949 <- mkDebugOperation(mod_1949_inner, "mod_1949");
    Operation_IFC mod_1950_inner <- mkFlatten(0);
    Operation_IFC mod_1950 <- mkDebugOperation(mod_1950_inner, "mod_1950");
    Operation_IFC mod_1951_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1951 <- mkDebugOperation(mod_1951_inner, "mod_1951");
    Operation_IFC mod_1952_inner <- mkUnaryMap(1749, silu_tile);
    Operation_IFC mod_1952 <- mkDebugOperation(mod_1952_inner, "mod_1952");
    Operation_IFC mod_1953_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1953 <- mkDebugOperation(mod_1953_inner, "mod_1953");
    Operation_IFC mod_1954_inner <- mkBinaryMap(1621, matmul_t_tile);
    Operation_IFC mod_1954 <- mkDebugOperation(mod_1954_inner, "mod_1954");
    PMU_IFC mod_1955_bufferize <- mkPMU(2);
    Operation_IFC mod_1955_inner = mod_1955_bufferize.operation;
    Operation_IFC mod_1955 <- mkDebugOperation(mod_1955_inner, "mod_1955");
    Operation_IFC mod_1956_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1956 <- mkDebugOperation(mod_1956_inner, "mod_1956");
    Operation_IFC mod_1957_inner <- mkFlatten(1);
    Operation_IFC mod_1957 <- mkDebugOperation(mod_1957_inner, "mod_1957");
    Operation_IFC mod_1958_inner <- mkFlatten(0);
    Operation_IFC mod_1958 <- mkDebugOperation(mod_1958_inner, "mod_1958");
    PMU_IFC mod_1959_bufferize <- mkPMU(1);
    Operation_IFC mod_1959_inner = mod_1959_bufferize.operation;
    Operation_IFC mod_1959 <- mkDebugOperation(mod_1959_inner, "mod_1959");
    Operation_IFC mod_1960_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1960 <- mkDebugOperation(mod_1960_inner, "mod_1960");
    PMU_IFC mod_1961_bufferize <- mkPMU(2);
    Operation_IFC mod_1961_inner = mod_1961_bufferize.operation;
    Operation_IFC mod_1961 <- mkDebugOperation(mod_1961_inner, "mod_1961");
    Operation_IFC mod_1962_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1962 <- mkDebugOperation(mod_1962_inner, "mod_1962");
    Operation_IFC mod_1963_inner <- mkFlatten(1);
    Operation_IFC mod_1963 <- mkDebugOperation(mod_1963_inner, "mod_1963");
    Operation_IFC mod_1964_inner <- mkFlatten(0);
    Operation_IFC mod_1964 <- mkDebugOperation(mod_1964_inner, "mod_1964");
    Operation_IFC mod_1965_inner <- mkRepeatStatic(16);
    Operation_IFC mod_1965 <- mkDebugOperation(mod_1965_inner, "mod_1965");
    Operation_IFC mod_1966_inner <- mkRepeatStatic(2);
    Operation_IFC mod_1966 <- mkDebugOperation(mod_1966_inner, "mod_1966");
    PMU_IFC mod_1967_bufferize <- mkPMU(2);
    Operation_IFC mod_1967_inner = mod_1967_bufferize.operation;
    Operation_IFC mod_1967 <- mkDebugOperation(mod_1967_inner, "mod_1967");
    rule rule_2492;
        ChannelMessage t;
        t <- mod_1941.get(0);
        mod_1942.put(0, t);
    endrule
    rule rule_2493;
        ChannelMessage t;
        t <- mod_1940.get(0);
        mod_1941.put(0, t);
    endrule
    rule rule_2494;
        ChannelMessage t;
        t <- mod_1963.get(0);
        mod_1961.put(0, t);
    endrule
    rule rule_2495;
        ChannelMessage t;
        t <- mod_1964.get(0);
        mod_1963.put(0, t);
    endrule
    rule rule_2496;
        ChannelMessage t;
        t <- mod_1948.get(0);
        mod_1947.put(1, t);
    endrule
    rule rule_2497;
        ChannelMessage t;
        t <- mod_1931.get(0);
        mod_1967.put(0, t);
    endrule
    rule rule_2498;
        ChannelMessage t;
        t <- mod_1947.get(0);
        mod_1948.put(0, t);
    endrule
    rule rule_2499;
        ChannelMessage t;
        t <- mod_1946.get(0);
        mod_1946.put(1, t);
    endrule
    rule rule_2500;
        ChannelMessage t;
        t <- mod_1960.get(0);
        mod_1959.put(1, t);
    endrule
    rule rule_2501;
        ChannelMessage t;
        t <- mod_1952.get(0);
        mod_1938.put(1, t);
    endrule
    rule rule_2502;
        ChannelMessage t;
        t <- mod_1939.get(1);
        mod_1940.put(0, t);
    endrule
    rule rule_2503;
        ChannelMessage t;
        t <- mod_1966.get(0);
        mod_1933.put(1, t);
    endrule
    rule rule_2504;
        ChannelMessage t;
        t <- mod_1958.get(0);
        mod_1957.put(0, t);
    endrule
    rule rule_2505;
        ChannelMessage t;
        t <- mod_1953.get(0);
        mod_1952.put(0, t);
    endrule
    rule rule_2506;
        ChannelMessage t;
        t <- mod_1967.get(0);
        mod_1967.put(1, t);
    endrule
    rule rule_2507;
        ChannelMessage t;
        t <- mod_1967.get(1);
        mod_1931.put(1, t);
    endrule
    rule rule_2508;
        ChannelMessage t;
        t <- mod_1965.get(0);
        mod_1935.put(1, t);
    endrule
    rule rule_2509;
        ChannelMessage t;
        t <- mod_1946.get(1);
        mod_1942.put(1, t);
    endrule
    rule rule_2510;
        ChannelMessage t;
        t <- mod_1961.get(1);
        mod_1936.put(1, t);
    endrule
    rule rule_2511;
        ChannelMessage t;
        t <- mod_1930.get(0);
        mod_1931.put(0, t);
    endrule
    rule rule_2512;
        ChannelMessage t;
        t <- mod_1959.get(0);
        mod_1960.put(0, t);
    endrule
    rule rule_2513;
        ChannelMessage t;
        t <- mod_1942.get(1);
        mod_1943.put(0, t);
    endrule
    rule rule_2514;
        ChannelMessage t;
        t <- mod_1936.get(0);
        mod_1937.put(0, t);
    endrule
    rule rule_2515;
        ChannelMessage t;
        t <- mod_1962.get(0);
        mod_1961.put(1, t);
    endrule
    rule rule_2516;
        ChannelMessage t;
        t <- mod_1934.get(0);
        mod_1959.put(0, t);
    endrule
    rule rule_2517;
        ChannelMessage t;
        t <- mod_1945.get(0);
        mod_1945.put(1, t);
    endrule
    rule rule_2518;
        ChannelMessage t;
        t <- mod_1928.get(0);
        mod_1929.put(0, t);
    endrule
    rule rule_2519;
        ChannelMessage t;
        t <- mod_1939.get(0);
        mod_1951.put(0, t);
    endrule
    rule rule_2520;
        ChannelMessage t;
        t <- mod_1943.get(0);
        mod_1945.put(0, t);
    endrule
    rule rule_2521;
        ChannelMessage t;
        t <- mod_1937.get(0);
        mod_1938.put(0, t);
    endrule
    rule rule_2522;
        ChannelMessage t;
        t <- mod_1933.get(1);
        mod_1934.put(0, t);
    endrule
    rule rule_2523;
        ChannelMessage t;
        t <- mod_1951.get(0);
        mod_1939.put(1, t);
    endrule
    rule rule_2524;
        ChannelMessage t;
        t <- mod_1932.get(3);
        mod_1933.put(0, t);
    endrule
    rule rule_2525;
        ChannelMessage t;
        t <- mod_1943.get(1);
        mod_1944.put(1, t);
    endrule
    rule rule_2526;
        ChannelMessage t;
        t <- mod_1954.get(0);
        mod_1953.put(0, t);
    endrule
    rule rule_2527;
        ChannelMessage t;
        t <- mod_1942.get(0);
        mod_1946.put(0, t);
    endrule
    rule rule_2528;
        ChannelMessage t;
        t <- mod_1959.get(1);
        mod_1954.put(0, t);
    endrule
    rule rule_2529;
        ChannelMessage t;
        t <- mod_1933.get(0);
        mod_1966.put(0, t);
    endrule
    rule rule_2530;
        ChannelMessage t;
        t <- mod_1929.get(0);
        mod_1930.put(0, t);
    endrule
    rule rule_2531;
        ChannelMessage t;
        t <- mod_1950.get(0);
        mod_1949.put(0, t);
    endrule
    rule rule_2532;
        ChannelMessage t;
        t <- mod_1955.get(0);
        mod_1956.put(0, t);
    endrule
    rule rule_2533;
        ChannelMessage t;
        t <- mod_1947.get(1);
        mod_1940.put(1, t);
    endrule
    rule rule_2534;
        ChannelMessage t;
        t <- mod_1935.get(0);
        mod_1965.put(0, t);
    endrule
    rule rule_2535;
        ChannelMessage t;
        t <- mod_1949.get(0);
        mod_1947.put(0, t);
    endrule
    rule rule_2536;
        ChannelMessage t;
        t <- mod_1934.get(1);
        mod_1935.put(0, t);
    endrule
    rule rule_2537;
        ChannelMessage t;
        t <- mod_1961.get(0);
        mod_1962.put(0, t);
    endrule
    rule rule_2538;
        ChannelMessage t;
        t <- mod_1931.get(1);
        mod_1932.put(0, t);
    endrule
    rule rule_2539;
        ChannelMessage t;
        t <- mod_1956.get(0);
        mod_1955.put(1, t);
    endrule
    rule rule_2540;
        ChannelMessage t;
        t <- mod_1938.get(0);
        mod_1939.put(0, t);
    endrule
    rule rule_2541;
        ChannelMessage t;
        t <- mod_1945.get(1);
        mod_1943.put(1, t);
    endrule
    rule rule_2542;
        ChannelMessage t;
        t <- mod_1955.get(1);
        mod_1954.put(1, t);
    endrule
    rule rule_2543;
        ChannelMessage t;
        t <- mod_1957.get(0);
        mod_1955.put(0, t);
    endrule
    rule rule_2544;
        ChannelMessage t;
        t <- mod_1935.get(1);
        mod_1936.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1928.put(0, t);
        end
        if (i == 1) begin
            mod_1944.put(0, t);
        end
        if (i == 2) begin
            mod_1950.put(0, t);
        end
        if (i == 3) begin
            mod_1958.put(0, t);
        end
        if (i == 4) begin
            mod_1964.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 2) begin
            t <- mod_1932.get(0);
        end
        if (i == 0) begin
            t <- mod_1932.get(1);
        end
        if (i == 3) begin
            t <- mod_1932.get(2);
        end
        if (i == 1) begin
            t <- mod_1944.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6082 (Operation_IFC);
    Operation_IFC mod_1969_inner <- mkReshape(2, 64);
    Operation_IFC mod_1969 <- mkDebugOperation(mod_1969_inner, "mod_1969");
    Operation_IFC mod_1970_inner <- mkFlatten(1);
    Operation_IFC mod_1970 <- mkDebugOperation(mod_1970_inner, "mod_1970");
    Operation_IFC mod_1971_inner <- mkFlatten(2);
    Operation_IFC mod_1971 <- mkDebugOperation(mod_1971_inner, "mod_1971");
    Operation_IFC mod_1972_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_1972 <- mkDebugOperation(mod_1972_inner, "mod_1972");
    Broadcast_IFC#(4) mod_1973_inner <- mkBroadcast(4);
    Operation_IFC mod_1973 <- mkDebugOperation(mod_1973_inner.op, "mod_1973");
    PMU_IFC mod_1974_bufferize <- mkPMU(2);
    Operation_IFC mod_1974_inner = mod_1974_bufferize.operation;
    Operation_IFC mod_1974 <- mkDebugOperation(mod_1974_inner, "mod_1974");
    Broadcast_IFC#(2) mod_1975_inner <- mkBroadcast(2);
    Operation_IFC mod_1975 <- mkDebugOperation(mod_1975_inner.op, "mod_1975");
    PMU_IFC mod_1976_bufferize <- mkPMU(1);
    Operation_IFC mod_1976_inner = mod_1976_bufferize.operation;
    Operation_IFC mod_1976 <- mkDebugOperation(mod_1976_inner, "mod_1976");
    Operation_IFC mod_1977_inner <- mkBinaryMap(1108, matmul_t_tile);
    Operation_IFC mod_1977 <- mkDebugOperation(mod_1977_inner, "mod_1977");
    Operation_IFC mod_1978_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1978 <- mkDebugOperation(mod_1978_inner, "mod_1978");
    Operation_IFC mod_1979_inner <- mkBinaryMap(1876, mul_tile);
    Operation_IFC mod_1979 <- mkDebugOperation(mod_1979_inner, "mod_1979");
    PMU_IFC mod_1980_bufferize <- mkPMU(1);
    Operation_IFC mod_1980_inner = mod_1980_bufferize.operation;
    Operation_IFC mod_1980 <- mkDebugOperation(mod_1980_inner, "mod_1980");
    Operation_IFC mod_1981_inner <- mkBinaryMap(2467, matmul_t_tile);
    Operation_IFC mod_1981 <- mkDebugOperation(mod_1981_inner, "mod_1981");
    Operation_IFC mod_1982_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1982 <- mkDebugOperation(mod_1982_inner, "mod_1982");
    Operation_IFC mod_1983_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_1983 <- mkDebugOperation(mod_1983_inner, "mod_1983");
    Operation_IFC mod_1984_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_1984 <- mkDebugOperation(mod_1984_inner, "mod_1984");
    Operation_IFC mod_1985_inner <- mkBinaryMap(2775, mul_tile);
    Operation_IFC mod_1985 <- mkDebugOperation(mod_1985_inner, "mod_1985");
    PMU_IFC mod_1986_bufferize <- mkPMU(1);
    Operation_IFC mod_1986_inner = mod_1986_bufferize.operation;
    Operation_IFC mod_1986 <- mkDebugOperation(mod_1986_inner, "mod_1986");
    PMU_IFC mod_1987_bufferize <- mkPMU(2);
    Operation_IFC mod_1987_inner = mod_1987_bufferize.operation;
    Operation_IFC mod_1987 <- mkDebugOperation(mod_1987_inner, "mod_1987");
    PMU_IFC mod_1988_bufferize <- mkPMU(2);
    Operation_IFC mod_1988_inner = mod_1988_bufferize.operation;
    Operation_IFC mod_1988 <- mkDebugOperation(mod_1988_inner, "mod_1988");
    Operation_IFC mod_1989_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1989 <- mkDebugOperation(mod_1989_inner, "mod_1989");
    Operation_IFC mod_1990_inner <- mkFlatten(1);
    Operation_IFC mod_1990 <- mkDebugOperation(mod_1990_inner, "mod_1990");
    Operation_IFC mod_1991_inner <- mkFlatten(0);
    Operation_IFC mod_1991 <- mkDebugOperation(mod_1991_inner, "mod_1991");
    Operation_IFC mod_1992_inner <- mkRepeatStatic(3);
    Operation_IFC mod_1992 <- mkDebugOperation(mod_1992_inner, "mod_1992");
    Operation_IFC mod_1993_inner <- mkUnaryMap(1748, silu_tile);
    Operation_IFC mod_1993 <- mkDebugOperation(mod_1993_inner, "mod_1993");
    Operation_IFC mod_1994_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_1994 <- mkDebugOperation(mod_1994_inner, "mod_1994");
    Operation_IFC mod_1995_inner <- mkBinaryMap(1620, matmul_t_tile);
    Operation_IFC mod_1995 <- mkDebugOperation(mod_1995_inner, "mod_1995");
    PMU_IFC mod_1996_bufferize <- mkPMU(2);
    Operation_IFC mod_1996_inner = mod_1996_bufferize.operation;
    Operation_IFC mod_1996 <- mkDebugOperation(mod_1996_inner, "mod_1996");
    Operation_IFC mod_1997_inner <- mkRepeatStatic(8);
    Operation_IFC mod_1997 <- mkDebugOperation(mod_1997_inner, "mod_1997");
    Operation_IFC mod_1998_inner <- mkFlatten(1);
    Operation_IFC mod_1998 <- mkDebugOperation(mod_1998_inner, "mod_1998");
    Operation_IFC mod_1999_inner <- mkFlatten(0);
    Operation_IFC mod_1999 <- mkDebugOperation(mod_1999_inner, "mod_1999");
    PMU_IFC mod_2000_bufferize <- mkPMU(1);
    Operation_IFC mod_2000_inner = mod_2000_bufferize.operation;
    Operation_IFC mod_2000 <- mkDebugOperation(mod_2000_inner, "mod_2000");
    Operation_IFC mod_2001_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2001 <- mkDebugOperation(mod_2001_inner, "mod_2001");
    PMU_IFC mod_2002_bufferize <- mkPMU(2);
    Operation_IFC mod_2002_inner = mod_2002_bufferize.operation;
    Operation_IFC mod_2002 <- mkDebugOperation(mod_2002_inner, "mod_2002");
    Operation_IFC mod_2003_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2003 <- mkDebugOperation(mod_2003_inner, "mod_2003");
    Operation_IFC mod_2004_inner <- mkFlatten(1);
    Operation_IFC mod_2004 <- mkDebugOperation(mod_2004_inner, "mod_2004");
    Operation_IFC mod_2005_inner <- mkFlatten(0);
    Operation_IFC mod_2005 <- mkDebugOperation(mod_2005_inner, "mod_2005");
    Operation_IFC mod_2006_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2006 <- mkDebugOperation(mod_2006_inner, "mod_2006");
    Operation_IFC mod_2007_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2007 <- mkDebugOperation(mod_2007_inner, "mod_2007");
    PMU_IFC mod_2008_bufferize <- mkPMU(2);
    Operation_IFC mod_2008_inner = mod_2008_bufferize.operation;
    Operation_IFC mod_2008 <- mkDebugOperation(mod_2008_inner, "mod_2008");
    rule rule_2545;
        ChannelMessage t;
        t <- mod_1994.get(0);
        mod_1993.put(0, t);
    endrule
    rule rule_2546;
        ChannelMessage t;
        t <- mod_1971.get(0);
        mod_1972.put(0, t);
    endrule
    rule rule_2547;
        ChannelMessage t;
        t <- mod_2003.get(0);
        mod_2002.put(1, t);
    endrule
    rule rule_2548;
        ChannelMessage t;
        t <- mod_1984.get(0);
        mod_1986.put(0, t);
    endrule
    rule rule_2549;
        ChannelMessage t;
        t <- mod_1979.get(0);
        mod_1980.put(0, t);
    endrule
    rule rule_2550;
        ChannelMessage t;
        t <- mod_1970.get(0);
        mod_1971.put(0, t);
    endrule
    rule rule_2551;
        ChannelMessage t;
        t <- mod_1996.get(1);
        mod_1995.put(1, t);
    endrule
    rule rule_2552;
        ChannelMessage t;
        t <- mod_1983.get(0);
        mod_1987.put(0, t);
    endrule
    rule rule_2553;
        ChannelMessage t;
        t <- mod_1988.get(1);
        mod_1981.put(1, t);
    endrule
    rule rule_2554;
        ChannelMessage t;
        t <- mod_2000.get(0);
        mod_2001.put(0, t);
    endrule
    rule rule_2555;
        ChannelMessage t;
        t <- mod_2008.get(1);
        mod_1972.put(1, t);
    endrule
    rule rule_2556;
        ChannelMessage t;
        t <- mod_1980.get(1);
        mod_1981.put(0, t);
    endrule
    rule rule_2557;
        ChannelMessage t;
        t <- mod_2000.get(1);
        mod_1995.put(0, t);
    endrule
    rule rule_2558;
        ChannelMessage t;
        t <- mod_1982.get(0);
        mod_1983.put(0, t);
    endrule
    rule rule_2559;
        ChannelMessage t;
        t <- mod_2008.get(0);
        mod_2008.put(1, t);
    endrule
    rule rule_2560;
        ChannelMessage t;
        t <- mod_2004.get(0);
        mod_2002.put(0, t);
    endrule
    rule rule_2561;
        ChannelMessage t;
        t <- mod_1999.get(0);
        mod_1998.put(0, t);
    endrule
    rule rule_2562;
        ChannelMessage t;
        t <- mod_1987.get(0);
        mod_1987.put(1, t);
    endrule
    rule rule_2563;
        ChannelMessage t;
        t <- mod_1992.get(0);
        mod_1980.put(1, t);
    endrule
    rule rule_2564;
        ChannelMessage t;
        t <- mod_1988.get(0);
        mod_1989.put(0, t);
    endrule
    rule rule_2565;
        ChannelMessage t;
        t <- mod_1996.get(0);
        mod_1997.put(0, t);
    endrule
    rule rule_2566;
        ChannelMessage t;
        t <- mod_2001.get(0);
        mod_2000.put(1, t);
    endrule
    rule rule_2567;
        ChannelMessage t;
        t <- mod_1998.get(0);
        mod_1996.put(0, t);
    endrule
    rule rule_2568;
        ChannelMessage t;
        t <- mod_1977.get(0);
        mod_1978.put(0, t);
    endrule
    rule rule_2569;
        ChannelMessage t;
        t <- mod_1978.get(0);
        mod_1979.put(0, t);
    endrule
    rule rule_2570;
        ChannelMessage t;
        t <- mod_1972.get(1);
        mod_1973.put(0, t);
    endrule
    rule rule_2571;
        ChannelMessage t;
        t <- mod_2007.get(0);
        mod_1974.put(1, t);
    endrule
    rule rule_2572;
        ChannelMessage t;
        t <- mod_1991.get(0);
        mod_1990.put(0, t);
    endrule
    rule rule_2573;
        ChannelMessage t;
        t <- mod_1986.get(0);
        mod_1986.put(1, t);
    endrule
    rule rule_2574;
        ChannelMessage t;
        t <- mod_1976.get(1);
        mod_1977.put(0, t);
    endrule
    rule rule_2575;
        ChannelMessage t;
        t <- mod_1969.get(0);
        mod_1970.put(0, t);
    endrule
    rule rule_2576;
        ChannelMessage t;
        t <- mod_1986.get(1);
        mod_1984.put(1, t);
    endrule
    rule rule_2577;
        ChannelMessage t;
        t <- mod_1995.get(0);
        mod_1994.put(0, t);
    endrule
    rule rule_2578;
        ChannelMessage t;
        t <- mod_1973.get(3);
        mod_1974.put(0, t);
    endrule
    rule rule_2579;
        ChannelMessage t;
        t <- mod_1976.get(0);
        mod_2006.put(0, t);
    endrule
    rule rule_2580;
        ChannelMessage t;
        t <- mod_1997.get(0);
        mod_1996.put(1, t);
    endrule
    rule rule_2581;
        ChannelMessage t;
        t <- mod_1987.get(1);
        mod_1983.put(1, t);
    endrule
    rule rule_2582;
        ChannelMessage t;
        t <- mod_1972.get(0);
        mod_2008.put(0, t);
    endrule
    rule rule_2583;
        ChannelMessage t;
        t <- mod_1974.get(1);
        mod_1975.put(0, t);
    endrule
    rule rule_2584;
        ChannelMessage t;
        t <- mod_1990.get(0);
        mod_1988.put(0, t);
    endrule
    rule rule_2585;
        ChannelMessage t;
        t <- mod_1989.get(0);
        mod_1988.put(1, t);
    endrule
    rule rule_2586;
        ChannelMessage t;
        t <- mod_1974.get(0);
        mod_2007.put(0, t);
    endrule
    rule rule_2587;
        ChannelMessage t;
        t <- mod_2006.get(0);
        mod_1976.put(1, t);
    endrule
    rule rule_2588;
        ChannelMessage t;
        t <- mod_1984.get(1);
        mod_1985.put(1, t);
    endrule
    rule rule_2589;
        ChannelMessage t;
        t <- mod_1975.get(1);
        mod_1976.put(0, t);
    endrule
    rule rule_2590;
        ChannelMessage t;
        t <- mod_1981.get(0);
        mod_1982.put(0, t);
    endrule
    rule rule_2591;
        ChannelMessage t;
        t <- mod_1983.get(1);
        mod_1984.put(0, t);
    endrule
    rule rule_2592;
        ChannelMessage t;
        t <- mod_2002.get(1);
        mod_1977.put(1, t);
    endrule
    rule rule_2593;
        ChannelMessage t;
        t <- mod_1975.get(0);
        mod_2000.put(0, t);
    endrule
    rule rule_2594;
        ChannelMessage t;
        t <- mod_2002.get(0);
        mod_2003.put(0, t);
    endrule
    rule rule_2595;
        ChannelMessage t;
        t <- mod_2005.get(0);
        mod_2004.put(0, t);
    endrule
    rule rule_2596;
        ChannelMessage t;
        t <- mod_1993.get(0);
        mod_1979.put(1, t);
    endrule
    rule rule_2597;
        ChannelMessage t;
        t <- mod_1980.get(0);
        mod_1992.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1969.put(0, t);
        end
        if (i == 1) begin
            mod_1985.put(0, t);
        end
        if (i == 2) begin
            mod_1991.put(0, t);
        end
        if (i == 3) begin
            mod_1999.put(0, t);
        end
        if (i == 4) begin
            mod_2005.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_1973.get(0);
        end
        if (i == 1) begin
            t <- mod_1973.get(1);
        end
        if (i == 3) begin
            t <- mod_1973.get(2);
        end
        if (i == 2) begin
            t <- mod_1985.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6083 (Operation_IFC);
    Operation_IFC mod_2010_inner <- mkReshape(2, 64);
    Operation_IFC mod_2010 <- mkDebugOperation(mod_2010_inner, "mod_2010");
    Operation_IFC mod_2011_inner <- mkFlatten(1);
    Operation_IFC mod_2011 <- mkDebugOperation(mod_2011_inner, "mod_2011");
    Operation_IFC mod_2012_inner <- mkFlatten(2);
    Operation_IFC mod_2012 <- mkDebugOperation(mod_2012_inner, "mod_2012");
    Operation_IFC mod_2013_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2013 <- mkDebugOperation(mod_2013_inner, "mod_2013");
    Broadcast_IFC#(4) mod_2014_inner <- mkBroadcast(4);
    Operation_IFC mod_2014 <- mkDebugOperation(mod_2014_inner.op, "mod_2014");
    PMU_IFC mod_2015_bufferize <- mkPMU(2);
    Operation_IFC mod_2015_inner = mod_2015_bufferize.operation;
    Operation_IFC mod_2015 <- mkDebugOperation(mod_2015_inner, "mod_2015");
    Broadcast_IFC#(2) mod_2016_inner <- mkBroadcast(2);
    Operation_IFC mod_2016 <- mkDebugOperation(mod_2016_inner.op, "mod_2016");
    PMU_IFC mod_2017_bufferize <- mkPMU(1);
    Operation_IFC mod_2017_inner = mod_2017_bufferize.operation;
    Operation_IFC mod_2017 <- mkDebugOperation(mod_2017_inner, "mod_2017");
    Operation_IFC mod_2018_inner <- mkBinaryMap(1107, matmul_t_tile);
    Operation_IFC mod_2018 <- mkDebugOperation(mod_2018_inner, "mod_2018");
    Operation_IFC mod_2019_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2019 <- mkDebugOperation(mod_2019_inner, "mod_2019");
    Operation_IFC mod_2020_inner <- mkBinaryMap(1875, mul_tile);
    Operation_IFC mod_2020 <- mkDebugOperation(mod_2020_inner, "mod_2020");
    PMU_IFC mod_2021_bufferize <- mkPMU(1);
    Operation_IFC mod_2021_inner = mod_2021_bufferize.operation;
    Operation_IFC mod_2021 <- mkDebugOperation(mod_2021_inner, "mod_2021");
    Operation_IFC mod_2022_inner <- mkBinaryMap(2465, matmul_t_tile);
    Operation_IFC mod_2022 <- mkDebugOperation(mod_2022_inner, "mod_2022");
    Operation_IFC mod_2023_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2023 <- mkDebugOperation(mod_2023_inner, "mod_2023");
    Operation_IFC mod_2024_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2024 <- mkDebugOperation(mod_2024_inner, "mod_2024");
    Operation_IFC mod_2025_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2025 <- mkDebugOperation(mod_2025_inner, "mod_2025");
    Operation_IFC mod_2026_inner <- mkBinaryMap(2774, mul_tile);
    Operation_IFC mod_2026 <- mkDebugOperation(mod_2026_inner, "mod_2026");
    PMU_IFC mod_2027_bufferize <- mkPMU(1);
    Operation_IFC mod_2027_inner = mod_2027_bufferize.operation;
    Operation_IFC mod_2027 <- mkDebugOperation(mod_2027_inner, "mod_2027");
    PMU_IFC mod_2028_bufferize <- mkPMU(2);
    Operation_IFC mod_2028_inner = mod_2028_bufferize.operation;
    Operation_IFC mod_2028 <- mkDebugOperation(mod_2028_inner, "mod_2028");
    PMU_IFC mod_2029_bufferize <- mkPMU(2);
    Operation_IFC mod_2029_inner = mod_2029_bufferize.operation;
    Operation_IFC mod_2029 <- mkDebugOperation(mod_2029_inner, "mod_2029");
    Operation_IFC mod_2030_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2030 <- mkDebugOperation(mod_2030_inner, "mod_2030");
    Operation_IFC mod_2031_inner <- mkFlatten(1);
    Operation_IFC mod_2031 <- mkDebugOperation(mod_2031_inner, "mod_2031");
    Operation_IFC mod_2032_inner <- mkFlatten(0);
    Operation_IFC mod_2032 <- mkDebugOperation(mod_2032_inner, "mod_2032");
    Operation_IFC mod_2033_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2033 <- mkDebugOperation(mod_2033_inner, "mod_2033");
    Operation_IFC mod_2034_inner <- mkUnaryMap(1747, silu_tile);
    Operation_IFC mod_2034 <- mkDebugOperation(mod_2034_inner, "mod_2034");
    Operation_IFC mod_2035_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2035 <- mkDebugOperation(mod_2035_inner, "mod_2035");
    Operation_IFC mod_2036_inner <- mkBinaryMap(1619, matmul_t_tile);
    Operation_IFC mod_2036 <- mkDebugOperation(mod_2036_inner, "mod_2036");
    PMU_IFC mod_2037_bufferize <- mkPMU(2);
    Operation_IFC mod_2037_inner = mod_2037_bufferize.operation;
    Operation_IFC mod_2037 <- mkDebugOperation(mod_2037_inner, "mod_2037");
    Operation_IFC mod_2038_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2038 <- mkDebugOperation(mod_2038_inner, "mod_2038");
    Operation_IFC mod_2039_inner <- mkFlatten(1);
    Operation_IFC mod_2039 <- mkDebugOperation(mod_2039_inner, "mod_2039");
    Operation_IFC mod_2040_inner <- mkFlatten(0);
    Operation_IFC mod_2040 <- mkDebugOperation(mod_2040_inner, "mod_2040");
    PMU_IFC mod_2041_bufferize <- mkPMU(1);
    Operation_IFC mod_2041_inner = mod_2041_bufferize.operation;
    Operation_IFC mod_2041 <- mkDebugOperation(mod_2041_inner, "mod_2041");
    Operation_IFC mod_2042_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2042 <- mkDebugOperation(mod_2042_inner, "mod_2042");
    PMU_IFC mod_2043_bufferize <- mkPMU(2);
    Operation_IFC mod_2043_inner = mod_2043_bufferize.operation;
    Operation_IFC mod_2043 <- mkDebugOperation(mod_2043_inner, "mod_2043");
    Operation_IFC mod_2044_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2044 <- mkDebugOperation(mod_2044_inner, "mod_2044");
    Operation_IFC mod_2045_inner <- mkFlatten(1);
    Operation_IFC mod_2045 <- mkDebugOperation(mod_2045_inner, "mod_2045");
    Operation_IFC mod_2046_inner <- mkFlatten(0);
    Operation_IFC mod_2046 <- mkDebugOperation(mod_2046_inner, "mod_2046");
    Operation_IFC mod_2047_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2047 <- mkDebugOperation(mod_2047_inner, "mod_2047");
    Operation_IFC mod_2048_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2048 <- mkDebugOperation(mod_2048_inner, "mod_2048");
    PMU_IFC mod_2049_bufferize <- mkPMU(2);
    Operation_IFC mod_2049_inner = mod_2049_bufferize.operation;
    Operation_IFC mod_2049 <- mkDebugOperation(mod_2049_inner, "mod_2049");
    rule rule_2598;
        ChannelMessage t;
        t <- mod_2034.get(0);
        mod_2020.put(1, t);
    endrule
    rule rule_2599;
        ChannelMessage t;
        t <- mod_2021.get(1);
        mod_2022.put(0, t);
    endrule
    rule rule_2600;
        ChannelMessage t;
        t <- mod_2027.get(1);
        mod_2025.put(1, t);
    endrule
    rule rule_2601;
        ChannelMessage t;
        t <- mod_2037.get(1);
        mod_2036.put(1, t);
    endrule
    rule rule_2602;
        ChannelMessage t;
        t <- mod_2038.get(0);
        mod_2037.put(1, t);
    endrule
    rule rule_2603;
        ChannelMessage t;
        t <- mod_2045.get(0);
        mod_2043.put(0, t);
    endrule
    rule rule_2604;
        ChannelMessage t;
        t <- mod_2041.get(0);
        mod_2042.put(0, t);
    endrule
    rule rule_2605;
        ChannelMessage t;
        t <- mod_2019.get(0);
        mod_2020.put(0, t);
    endrule
    rule rule_2606;
        ChannelMessage t;
        t <- mod_2028.get(1);
        mod_2024.put(1, t);
    endrule
    rule rule_2607;
        ChannelMessage t;
        t <- mod_2035.get(0);
        mod_2034.put(0, t);
    endrule
    rule rule_2608;
        ChannelMessage t;
        t <- mod_2025.get(1);
        mod_2026.put(1, t);
    endrule
    rule rule_2609;
        ChannelMessage t;
        t <- mod_2024.get(0);
        mod_2028.put(0, t);
    endrule
    rule rule_2610;
        ChannelMessage t;
        t <- mod_2029.get(1);
        mod_2022.put(1, t);
    endrule
    rule rule_2611;
        ChannelMessage t;
        t <- mod_2041.get(1);
        mod_2036.put(0, t);
    endrule
    rule rule_2612;
        ChannelMessage t;
        t <- mod_2010.get(0);
        mod_2011.put(0, t);
    endrule
    rule rule_2613;
        ChannelMessage t;
        t <- mod_2027.get(0);
        mod_2027.put(1, t);
    endrule
    rule rule_2614;
        ChannelMessage t;
        t <- mod_2049.get(0);
        mod_2049.put(1, t);
    endrule
    rule rule_2615;
        ChannelMessage t;
        t <- mod_2028.get(0);
        mod_2028.put(1, t);
    endrule
    rule rule_2616;
        ChannelMessage t;
        t <- mod_2024.get(1);
        mod_2025.put(0, t);
    endrule
    rule rule_2617;
        ChannelMessage t;
        t <- mod_2021.get(0);
        mod_2033.put(0, t);
    endrule
    rule rule_2618;
        ChannelMessage t;
        t <- mod_2037.get(0);
        mod_2038.put(0, t);
    endrule
    rule rule_2619;
        ChannelMessage t;
        t <- mod_2047.get(0);
        mod_2017.put(1, t);
    endrule
    rule rule_2620;
        ChannelMessage t;
        t <- mod_2014.get(3);
        mod_2015.put(0, t);
    endrule
    rule rule_2621;
        ChannelMessage t;
        t <- mod_2015.get(1);
        mod_2016.put(0, t);
    endrule
    rule rule_2622;
        ChannelMessage t;
        t <- mod_2020.get(0);
        mod_2021.put(0, t);
    endrule
    rule rule_2623;
        ChannelMessage t;
        t <- mod_2016.get(1);
        mod_2017.put(0, t);
    endrule
    rule rule_2624;
        ChannelMessage t;
        t <- mod_2018.get(0);
        mod_2019.put(0, t);
    endrule
    rule rule_2625;
        ChannelMessage t;
        t <- mod_2025.get(0);
        mod_2027.put(0, t);
    endrule
    rule rule_2626;
        ChannelMessage t;
        t <- mod_2029.get(0);
        mod_2030.put(0, t);
    endrule
    rule rule_2627;
        ChannelMessage t;
        t <- mod_2013.get(0);
        mod_2049.put(0, t);
    endrule
    rule rule_2628;
        ChannelMessage t;
        t <- mod_2023.get(0);
        mod_2024.put(0, t);
    endrule
    rule rule_2629;
        ChannelMessage t;
        t <- mod_2046.get(0);
        mod_2045.put(0, t);
    endrule
    rule rule_2630;
        ChannelMessage t;
        t <- mod_2043.get(1);
        mod_2018.put(1, t);
    endrule
    rule rule_2631;
        ChannelMessage t;
        t <- mod_2033.get(0);
        mod_2021.put(1, t);
    endrule
    rule rule_2632;
        ChannelMessage t;
        t <- mod_2044.get(0);
        mod_2043.put(1, t);
    endrule
    rule rule_2633;
        ChannelMessage t;
        t <- mod_2022.get(0);
        mod_2023.put(0, t);
    endrule
    rule rule_2634;
        ChannelMessage t;
        t <- mod_2017.get(0);
        mod_2047.put(0, t);
    endrule
    rule rule_2635;
        ChannelMessage t;
        t <- mod_2032.get(0);
        mod_2031.put(0, t);
    endrule
    rule rule_2636;
        ChannelMessage t;
        t <- mod_2039.get(0);
        mod_2037.put(0, t);
    endrule
    rule rule_2637;
        ChannelMessage t;
        t <- mod_2040.get(0);
        mod_2039.put(0, t);
    endrule
    rule rule_2638;
        ChannelMessage t;
        t <- mod_2042.get(0);
        mod_2041.put(1, t);
    endrule
    rule rule_2639;
        ChannelMessage t;
        t <- mod_2013.get(1);
        mod_2014.put(0, t);
    endrule
    rule rule_2640;
        ChannelMessage t;
        t <- mod_2048.get(0);
        mod_2015.put(1, t);
    endrule
    rule rule_2641;
        ChannelMessage t;
        t <- mod_2015.get(0);
        mod_2048.put(0, t);
    endrule
    rule rule_2642;
        ChannelMessage t;
        t <- mod_2043.get(0);
        mod_2044.put(0, t);
    endrule
    rule rule_2643;
        ChannelMessage t;
        t <- mod_2017.get(1);
        mod_2018.put(0, t);
    endrule
    rule rule_2644;
        ChannelMessage t;
        t <- mod_2031.get(0);
        mod_2029.put(0, t);
    endrule
    rule rule_2645;
        ChannelMessage t;
        t <- mod_2012.get(0);
        mod_2013.put(0, t);
    endrule
    rule rule_2646;
        ChannelMessage t;
        t <- mod_2016.get(0);
        mod_2041.put(0, t);
    endrule
    rule rule_2647;
        ChannelMessage t;
        t <- mod_2011.get(0);
        mod_2012.put(0, t);
    endrule
    rule rule_2648;
        ChannelMessage t;
        t <- mod_2036.get(0);
        mod_2035.put(0, t);
    endrule
    rule rule_2649;
        ChannelMessage t;
        t <- mod_2030.get(0);
        mod_2029.put(1, t);
    endrule
    rule rule_2650;
        ChannelMessage t;
        t <- mod_2049.get(1);
        mod_2013.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2010.put(0, t);
        end
        if (i == 1) begin
            mod_2026.put(0, t);
        end
        if (i == 2) begin
            mod_2032.put(0, t);
        end
        if (i == 3) begin
            mod_2040.put(0, t);
        end
        if (i == 4) begin
            mod_2046.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_2014.get(0);
        end
        if (i == 3) begin
            t <- mod_2014.get(1);
        end
        if (i == 2) begin
            t <- mod_2014.get(2);
        end
        if (i == 1) begin
            t <- mod_2026.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6084 (Operation_IFC);
    Operation_IFC mod_2051_inner <- mkReshape(2, 64);
    Operation_IFC mod_2051 <- mkDebugOperation(mod_2051_inner, "mod_2051");
    Operation_IFC mod_2052_inner <- mkFlatten(1);
    Operation_IFC mod_2052 <- mkDebugOperation(mod_2052_inner, "mod_2052");
    Operation_IFC mod_2053_inner <- mkFlatten(2);
    Operation_IFC mod_2053 <- mkDebugOperation(mod_2053_inner, "mod_2053");
    Operation_IFC mod_2054_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2054 <- mkDebugOperation(mod_2054_inner, "mod_2054");
    Broadcast_IFC#(4) mod_2055_inner <- mkBroadcast(4);
    Operation_IFC mod_2055 <- mkDebugOperation(mod_2055_inner.op, "mod_2055");
    PMU_IFC mod_2056_bufferize <- mkPMU(2);
    Operation_IFC mod_2056_inner = mod_2056_bufferize.operation;
    Operation_IFC mod_2056 <- mkDebugOperation(mod_2056_inner, "mod_2056");
    Broadcast_IFC#(2) mod_2057_inner <- mkBroadcast(2);
    Operation_IFC mod_2057 <- mkDebugOperation(mod_2057_inner.op, "mod_2057");
    PMU_IFC mod_2058_bufferize <- mkPMU(1);
    Operation_IFC mod_2058_inner = mod_2058_bufferize.operation;
    Operation_IFC mod_2058 <- mkDebugOperation(mod_2058_inner, "mod_2058");
    Operation_IFC mod_2059_inner <- mkBinaryMap(1106, matmul_t_tile);
    Operation_IFC mod_2059 <- mkDebugOperation(mod_2059_inner, "mod_2059");
    Operation_IFC mod_2060_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2060 <- mkDebugOperation(mod_2060_inner, "mod_2060");
    Operation_IFC mod_2061_inner <- mkBinaryMap(1874, mul_tile);
    Operation_IFC mod_2061 <- mkDebugOperation(mod_2061_inner, "mod_2061");
    PMU_IFC mod_2062_bufferize <- mkPMU(1);
    Operation_IFC mod_2062_inner = mod_2062_bufferize.operation;
    Operation_IFC mod_2062 <- mkDebugOperation(mod_2062_inner, "mod_2062");
    Operation_IFC mod_2063_inner <- mkBinaryMap(2463, matmul_t_tile);
    Operation_IFC mod_2063 <- mkDebugOperation(mod_2063_inner, "mod_2063");
    Operation_IFC mod_2064_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2064 <- mkDebugOperation(mod_2064_inner, "mod_2064");
    Operation_IFC mod_2065_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2065 <- mkDebugOperation(mod_2065_inner, "mod_2065");
    Operation_IFC mod_2066_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2066 <- mkDebugOperation(mod_2066_inner, "mod_2066");
    Operation_IFC mod_2067_inner <- mkBinaryMap(2773, mul_tile);
    Operation_IFC mod_2067 <- mkDebugOperation(mod_2067_inner, "mod_2067");
    PMU_IFC mod_2068_bufferize <- mkPMU(1);
    Operation_IFC mod_2068_inner = mod_2068_bufferize.operation;
    Operation_IFC mod_2068 <- mkDebugOperation(mod_2068_inner, "mod_2068");
    PMU_IFC mod_2069_bufferize <- mkPMU(2);
    Operation_IFC mod_2069_inner = mod_2069_bufferize.operation;
    Operation_IFC mod_2069 <- mkDebugOperation(mod_2069_inner, "mod_2069");
    PMU_IFC mod_2070_bufferize <- mkPMU(2);
    Operation_IFC mod_2070_inner = mod_2070_bufferize.operation;
    Operation_IFC mod_2070 <- mkDebugOperation(mod_2070_inner, "mod_2070");
    Operation_IFC mod_2071_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2071 <- mkDebugOperation(mod_2071_inner, "mod_2071");
    Operation_IFC mod_2072_inner <- mkFlatten(1);
    Operation_IFC mod_2072 <- mkDebugOperation(mod_2072_inner, "mod_2072");
    Operation_IFC mod_2073_inner <- mkFlatten(0);
    Operation_IFC mod_2073 <- mkDebugOperation(mod_2073_inner, "mod_2073");
    Operation_IFC mod_2074_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2074 <- mkDebugOperation(mod_2074_inner, "mod_2074");
    Operation_IFC mod_2075_inner <- mkUnaryMap(1746, silu_tile);
    Operation_IFC mod_2075 <- mkDebugOperation(mod_2075_inner, "mod_2075");
    Operation_IFC mod_2076_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2076 <- mkDebugOperation(mod_2076_inner, "mod_2076");
    Operation_IFC mod_2077_inner <- mkBinaryMap(1618, matmul_t_tile);
    Operation_IFC mod_2077 <- mkDebugOperation(mod_2077_inner, "mod_2077");
    PMU_IFC mod_2078_bufferize <- mkPMU(2);
    Operation_IFC mod_2078_inner = mod_2078_bufferize.operation;
    Operation_IFC mod_2078 <- mkDebugOperation(mod_2078_inner, "mod_2078");
    Operation_IFC mod_2079_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2079 <- mkDebugOperation(mod_2079_inner, "mod_2079");
    Operation_IFC mod_2080_inner <- mkFlatten(1);
    Operation_IFC mod_2080 <- mkDebugOperation(mod_2080_inner, "mod_2080");
    Operation_IFC mod_2081_inner <- mkFlatten(0);
    Operation_IFC mod_2081 <- mkDebugOperation(mod_2081_inner, "mod_2081");
    PMU_IFC mod_2082_bufferize <- mkPMU(1);
    Operation_IFC mod_2082_inner = mod_2082_bufferize.operation;
    Operation_IFC mod_2082 <- mkDebugOperation(mod_2082_inner, "mod_2082");
    Operation_IFC mod_2083_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2083 <- mkDebugOperation(mod_2083_inner, "mod_2083");
    PMU_IFC mod_2084_bufferize <- mkPMU(2);
    Operation_IFC mod_2084_inner = mod_2084_bufferize.operation;
    Operation_IFC mod_2084 <- mkDebugOperation(mod_2084_inner, "mod_2084");
    Operation_IFC mod_2085_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2085 <- mkDebugOperation(mod_2085_inner, "mod_2085");
    Operation_IFC mod_2086_inner <- mkFlatten(1);
    Operation_IFC mod_2086 <- mkDebugOperation(mod_2086_inner, "mod_2086");
    Operation_IFC mod_2087_inner <- mkFlatten(0);
    Operation_IFC mod_2087 <- mkDebugOperation(mod_2087_inner, "mod_2087");
    Operation_IFC mod_2088_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2088 <- mkDebugOperation(mod_2088_inner, "mod_2088");
    Operation_IFC mod_2089_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2089 <- mkDebugOperation(mod_2089_inner, "mod_2089");
    PMU_IFC mod_2090_bufferize <- mkPMU(2);
    Operation_IFC mod_2090_inner = mod_2090_bufferize.operation;
    Operation_IFC mod_2090 <- mkDebugOperation(mod_2090_inner, "mod_2090");
    rule rule_2651;
        ChannelMessage t;
        t <- mod_2058.get(1);
        mod_2059.put(0, t);
    endrule
    rule rule_2652;
        ChannelMessage t;
        t <- mod_2068.get(1);
        mod_2066.put(1, t);
    endrule
    rule rule_2653;
        ChannelMessage t;
        t <- mod_2070.get(1);
        mod_2063.put(1, t);
    endrule
    rule rule_2654;
        ChannelMessage t;
        t <- mod_2074.get(0);
        mod_2062.put(1, t);
    endrule
    rule rule_2655;
        ChannelMessage t;
        t <- mod_2089.get(0);
        mod_2056.put(1, t);
    endrule
    rule rule_2656;
        ChannelMessage t;
        t <- mod_2078.get(0);
        mod_2079.put(0, t);
    endrule
    rule rule_2657;
        ChannelMessage t;
        t <- mod_2071.get(0);
        mod_2070.put(1, t);
    endrule
    rule rule_2658;
        ChannelMessage t;
        t <- mod_2088.get(0);
        mod_2058.put(1, t);
    endrule
    rule rule_2659;
        ChannelMessage t;
        t <- mod_2076.get(0);
        mod_2075.put(0, t);
    endrule
    rule rule_2660;
        ChannelMessage t;
        t <- mod_2055.get(3);
        mod_2056.put(0, t);
    endrule
    rule rule_2661;
        ChannelMessage t;
        t <- mod_2052.get(0);
        mod_2053.put(0, t);
    endrule
    rule rule_2662;
        ChannelMessage t;
        t <- mod_2062.get(0);
        mod_2074.put(0, t);
    endrule
    rule rule_2663;
        ChannelMessage t;
        t <- mod_2051.get(0);
        mod_2052.put(0, t);
    endrule
    rule rule_2664;
        ChannelMessage t;
        t <- mod_2066.get(0);
        mod_2068.put(0, t);
    endrule
    rule rule_2665;
        ChannelMessage t;
        t <- mod_2078.get(1);
        mod_2077.put(1, t);
    endrule
    rule rule_2666;
        ChannelMessage t;
        t <- mod_2063.get(0);
        mod_2064.put(0, t);
    endrule
    rule rule_2667;
        ChannelMessage t;
        t <- mod_2064.get(0);
        mod_2065.put(0, t);
    endrule
    rule rule_2668;
        ChannelMessage t;
        t <- mod_2065.get(1);
        mod_2066.put(0, t);
    endrule
    rule rule_2669;
        ChannelMessage t;
        t <- mod_2054.get(0);
        mod_2090.put(0, t);
    endrule
    rule rule_2670;
        ChannelMessage t;
        t <- mod_2062.get(1);
        mod_2063.put(0, t);
    endrule
    rule rule_2671;
        ChannelMessage t;
        t <- mod_2082.get(1);
        mod_2077.put(0, t);
    endrule
    rule rule_2672;
        ChannelMessage t;
        t <- mod_2070.get(0);
        mod_2071.put(0, t);
    endrule
    rule rule_2673;
        ChannelMessage t;
        t <- mod_2090.get(1);
        mod_2054.put(1, t);
    endrule
    rule rule_2674;
        ChannelMessage t;
        t <- mod_2081.get(0);
        mod_2080.put(0, t);
    endrule
    rule rule_2675;
        ChannelMessage t;
        t <- mod_2065.get(0);
        mod_2069.put(0, t);
    endrule
    rule rule_2676;
        ChannelMessage t;
        t <- mod_2056.get(0);
        mod_2089.put(0, t);
    endrule
    rule rule_2677;
        ChannelMessage t;
        t <- mod_2087.get(0);
        mod_2086.put(0, t);
    endrule
    rule rule_2678;
        ChannelMessage t;
        t <- mod_2058.get(0);
        mod_2088.put(0, t);
    endrule
    rule rule_2679;
        ChannelMessage t;
        t <- mod_2073.get(0);
        mod_2072.put(0, t);
    endrule
    rule rule_2680;
        ChannelMessage t;
        t <- mod_2082.get(0);
        mod_2083.put(0, t);
    endrule
    rule rule_2681;
        ChannelMessage t;
        t <- mod_2056.get(1);
        mod_2057.put(0, t);
    endrule
    rule rule_2682;
        ChannelMessage t;
        t <- mod_2075.get(0);
        mod_2061.put(1, t);
    endrule
    rule rule_2683;
        ChannelMessage t;
        t <- mod_2079.get(0);
        mod_2078.put(1, t);
    endrule
    rule rule_2684;
        ChannelMessage t;
        t <- mod_2069.get(1);
        mod_2065.put(1, t);
    endrule
    rule rule_2685;
        ChannelMessage t;
        t <- mod_2086.get(0);
        mod_2084.put(0, t);
    endrule
    rule rule_2686;
        ChannelMessage t;
        t <- mod_2060.get(0);
        mod_2061.put(0, t);
    endrule
    rule rule_2687;
        ChannelMessage t;
        t <- mod_2072.get(0);
        mod_2070.put(0, t);
    endrule
    rule rule_2688;
        ChannelMessage t;
        t <- mod_2084.get(0);
        mod_2085.put(0, t);
    endrule
    rule rule_2689;
        ChannelMessage t;
        t <- mod_2057.get(1);
        mod_2058.put(0, t);
    endrule
    rule rule_2690;
        ChannelMessage t;
        t <- mod_2057.get(0);
        mod_2082.put(0, t);
    endrule
    rule rule_2691;
        ChannelMessage t;
        t <- mod_2059.get(0);
        mod_2060.put(0, t);
    endrule
    rule rule_2692;
        ChannelMessage t;
        t <- mod_2090.get(0);
        mod_2090.put(1, t);
    endrule
    rule rule_2693;
        ChannelMessage t;
        t <- mod_2085.get(0);
        mod_2084.put(1, t);
    endrule
    rule rule_2694;
        ChannelMessage t;
        t <- mod_2054.get(1);
        mod_2055.put(0, t);
    endrule
    rule rule_2695;
        ChannelMessage t;
        t <- mod_2066.get(1);
        mod_2067.put(1, t);
    endrule
    rule rule_2696;
        ChannelMessage t;
        t <- mod_2084.get(1);
        mod_2059.put(1, t);
    endrule
    rule rule_2697;
        ChannelMessage t;
        t <- mod_2061.get(0);
        mod_2062.put(0, t);
    endrule
    rule rule_2698;
        ChannelMessage t;
        t <- mod_2068.get(0);
        mod_2068.put(1, t);
    endrule
    rule rule_2699;
        ChannelMessage t;
        t <- mod_2053.get(0);
        mod_2054.put(0, t);
    endrule
    rule rule_2700;
        ChannelMessage t;
        t <- mod_2077.get(0);
        mod_2076.put(0, t);
    endrule
    rule rule_2701;
        ChannelMessage t;
        t <- mod_2069.get(0);
        mod_2069.put(1, t);
    endrule
    rule rule_2702;
        ChannelMessage t;
        t <- mod_2080.get(0);
        mod_2078.put(0, t);
    endrule
    rule rule_2703;
        ChannelMessage t;
        t <- mod_2083.get(0);
        mod_2082.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2051.put(0, t);
        end
        if (i == 1) begin
            mod_2067.put(0, t);
        end
        if (i == 2) begin
            mod_2073.put(0, t);
        end
        if (i == 3) begin
            mod_2081.put(0, t);
        end
        if (i == 4) begin
            mod_2087.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 2) begin
            t <- mod_2055.get(0);
        end
        if (i == 3) begin
            t <- mod_2055.get(1);
        end
        if (i == 1) begin
            t <- mod_2055.get(2);
        end
        if (i == 0) begin
            t <- mod_2067.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6085 (Operation_IFC);
    Operation_IFC mod_2092_inner <- mkReshape(2, 64);
    Operation_IFC mod_2092 <- mkDebugOperation(mod_2092_inner, "mod_2092");
    Operation_IFC mod_2093_inner <- mkFlatten(1);
    Operation_IFC mod_2093 <- mkDebugOperation(mod_2093_inner, "mod_2093");
    Operation_IFC mod_2094_inner <- mkFlatten(2);
    Operation_IFC mod_2094 <- mkDebugOperation(mod_2094_inner, "mod_2094");
    Operation_IFC mod_2095_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2095 <- mkDebugOperation(mod_2095_inner, "mod_2095");
    Broadcast_IFC#(4) mod_2096_inner <- mkBroadcast(4);
    Operation_IFC mod_2096 <- mkDebugOperation(mod_2096_inner.op, "mod_2096");
    PMU_IFC mod_2097_bufferize <- mkPMU(2);
    Operation_IFC mod_2097_inner = mod_2097_bufferize.operation;
    Operation_IFC mod_2097 <- mkDebugOperation(mod_2097_inner, "mod_2097");
    Broadcast_IFC#(2) mod_2098_inner <- mkBroadcast(2);
    Operation_IFC mod_2098 <- mkDebugOperation(mod_2098_inner.op, "mod_2098");
    PMU_IFC mod_2099_bufferize <- mkPMU(1);
    Operation_IFC mod_2099_inner = mod_2099_bufferize.operation;
    Operation_IFC mod_2099 <- mkDebugOperation(mod_2099_inner, "mod_2099");
    Operation_IFC mod_2100_inner <- mkBinaryMap(1105, matmul_t_tile);
    Operation_IFC mod_2100 <- mkDebugOperation(mod_2100_inner, "mod_2100");
    Operation_IFC mod_2101_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2101 <- mkDebugOperation(mod_2101_inner, "mod_2101");
    Operation_IFC mod_2102_inner <- mkBinaryMap(1873, mul_tile);
    Operation_IFC mod_2102 <- mkDebugOperation(mod_2102_inner, "mod_2102");
    PMU_IFC mod_2103_bufferize <- mkPMU(1);
    Operation_IFC mod_2103_inner = mod_2103_bufferize.operation;
    Operation_IFC mod_2103 <- mkDebugOperation(mod_2103_inner, "mod_2103");
    Operation_IFC mod_2104_inner <- mkBinaryMap(2461, matmul_t_tile);
    Operation_IFC mod_2104 <- mkDebugOperation(mod_2104_inner, "mod_2104");
    Operation_IFC mod_2105_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2105 <- mkDebugOperation(mod_2105_inner, "mod_2105");
    Operation_IFC mod_2106_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2106 <- mkDebugOperation(mod_2106_inner, "mod_2106");
    Operation_IFC mod_2107_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2107 <- mkDebugOperation(mod_2107_inner, "mod_2107");
    Operation_IFC mod_2108_inner <- mkBinaryMap(2772, mul_tile);
    Operation_IFC mod_2108 <- mkDebugOperation(mod_2108_inner, "mod_2108");
    PMU_IFC mod_2109_bufferize <- mkPMU(1);
    Operation_IFC mod_2109_inner = mod_2109_bufferize.operation;
    Operation_IFC mod_2109 <- mkDebugOperation(mod_2109_inner, "mod_2109");
    PMU_IFC mod_2110_bufferize <- mkPMU(2);
    Operation_IFC mod_2110_inner = mod_2110_bufferize.operation;
    Operation_IFC mod_2110 <- mkDebugOperation(mod_2110_inner, "mod_2110");
    PMU_IFC mod_2111_bufferize <- mkPMU(2);
    Operation_IFC mod_2111_inner = mod_2111_bufferize.operation;
    Operation_IFC mod_2111 <- mkDebugOperation(mod_2111_inner, "mod_2111");
    Operation_IFC mod_2112_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2112 <- mkDebugOperation(mod_2112_inner, "mod_2112");
    Operation_IFC mod_2113_inner <- mkFlatten(1);
    Operation_IFC mod_2113 <- mkDebugOperation(mod_2113_inner, "mod_2113");
    Operation_IFC mod_2114_inner <- mkFlatten(0);
    Operation_IFC mod_2114 <- mkDebugOperation(mod_2114_inner, "mod_2114");
    Operation_IFC mod_2115_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2115 <- mkDebugOperation(mod_2115_inner, "mod_2115");
    Operation_IFC mod_2116_inner <- mkUnaryMap(1745, silu_tile);
    Operation_IFC mod_2116 <- mkDebugOperation(mod_2116_inner, "mod_2116");
    Operation_IFC mod_2117_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2117 <- mkDebugOperation(mod_2117_inner, "mod_2117");
    Operation_IFC mod_2118_inner <- mkBinaryMap(1617, matmul_t_tile);
    Operation_IFC mod_2118 <- mkDebugOperation(mod_2118_inner, "mod_2118");
    PMU_IFC mod_2119_bufferize <- mkPMU(2);
    Operation_IFC mod_2119_inner = mod_2119_bufferize.operation;
    Operation_IFC mod_2119 <- mkDebugOperation(mod_2119_inner, "mod_2119");
    Operation_IFC mod_2120_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2120 <- mkDebugOperation(mod_2120_inner, "mod_2120");
    Operation_IFC mod_2121_inner <- mkFlatten(1);
    Operation_IFC mod_2121 <- mkDebugOperation(mod_2121_inner, "mod_2121");
    Operation_IFC mod_2122_inner <- mkFlatten(0);
    Operation_IFC mod_2122 <- mkDebugOperation(mod_2122_inner, "mod_2122");
    PMU_IFC mod_2123_bufferize <- mkPMU(1);
    Operation_IFC mod_2123_inner = mod_2123_bufferize.operation;
    Operation_IFC mod_2123 <- mkDebugOperation(mod_2123_inner, "mod_2123");
    Operation_IFC mod_2124_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2124 <- mkDebugOperation(mod_2124_inner, "mod_2124");
    PMU_IFC mod_2125_bufferize <- mkPMU(2);
    Operation_IFC mod_2125_inner = mod_2125_bufferize.operation;
    Operation_IFC mod_2125 <- mkDebugOperation(mod_2125_inner, "mod_2125");
    Operation_IFC mod_2126_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2126 <- mkDebugOperation(mod_2126_inner, "mod_2126");
    Operation_IFC mod_2127_inner <- mkFlatten(1);
    Operation_IFC mod_2127 <- mkDebugOperation(mod_2127_inner, "mod_2127");
    Operation_IFC mod_2128_inner <- mkFlatten(0);
    Operation_IFC mod_2128 <- mkDebugOperation(mod_2128_inner, "mod_2128");
    Operation_IFC mod_2129_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2129 <- mkDebugOperation(mod_2129_inner, "mod_2129");
    Operation_IFC mod_2130_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2130 <- mkDebugOperation(mod_2130_inner, "mod_2130");
    PMU_IFC mod_2131_bufferize <- mkPMU(2);
    Operation_IFC mod_2131_inner = mod_2131_bufferize.operation;
    Operation_IFC mod_2131 <- mkDebugOperation(mod_2131_inner, "mod_2131");
    rule rule_2704;
        ChannelMessage t;
        t <- mod_2116.get(0);
        mod_2102.put(1, t);
    endrule
    rule rule_2705;
        ChannelMessage t;
        t <- mod_2092.get(0);
        mod_2093.put(0, t);
    endrule
    rule rule_2706;
        ChannelMessage t;
        t <- mod_2099.get(0);
        mod_2129.put(0, t);
    endrule
    rule rule_2707;
        ChannelMessage t;
        t <- mod_2109.get(1);
        mod_2107.put(1, t);
    endrule
    rule rule_2708;
        ChannelMessage t;
        t <- mod_2099.get(1);
        mod_2100.put(0, t);
    endrule
    rule rule_2709;
        ChannelMessage t;
        t <- mod_2111.get(1);
        mod_2104.put(1, t);
    endrule
    rule rule_2710;
        ChannelMessage t;
        t <- mod_2107.get(1);
        mod_2108.put(1, t);
    endrule
    rule rule_2711;
        ChannelMessage t;
        t <- mod_2119.get(1);
        mod_2118.put(1, t);
    endrule
    rule rule_2712;
        ChannelMessage t;
        t <- mod_2114.get(0);
        mod_2113.put(0, t);
    endrule
    rule rule_2713;
        ChannelMessage t;
        t <- mod_2098.get(0);
        mod_2123.put(0, t);
    endrule
    rule rule_2714;
        ChannelMessage t;
        t <- mod_2130.get(0);
        mod_2097.put(1, t);
    endrule
    rule rule_2715;
        ChannelMessage t;
        t <- mod_2126.get(0);
        mod_2125.put(1, t);
    endrule
    rule rule_2716;
        ChannelMessage t;
        t <- mod_2122.get(0);
        mod_2121.put(0, t);
    endrule
    rule rule_2717;
        ChannelMessage t;
        t <- mod_2121.get(0);
        mod_2119.put(0, t);
    endrule
    rule rule_2718;
        ChannelMessage t;
        t <- mod_2111.get(0);
        mod_2112.put(0, t);
    endrule
    rule rule_2719;
        ChannelMessage t;
        t <- mod_2112.get(0);
        mod_2111.put(1, t);
    endrule
    rule rule_2720;
        ChannelMessage t;
        t <- mod_2097.get(1);
        mod_2098.put(0, t);
    endrule
    rule rule_2721;
        ChannelMessage t;
        t <- mod_2124.get(0);
        mod_2123.put(1, t);
    endrule
    rule rule_2722;
        ChannelMessage t;
        t <- mod_2102.get(0);
        mod_2103.put(0, t);
    endrule
    rule rule_2723;
        ChannelMessage t;
        t <- mod_2129.get(0);
        mod_2099.put(1, t);
    endrule
    rule rule_2724;
        ChannelMessage t;
        t <- mod_2106.get(1);
        mod_2107.put(0, t);
    endrule
    rule rule_2725;
        ChannelMessage t;
        t <- mod_2106.get(0);
        mod_2110.put(0, t);
    endrule
    rule rule_2726;
        ChannelMessage t;
        t <- mod_2101.get(0);
        mod_2102.put(0, t);
    endrule
    rule rule_2727;
        ChannelMessage t;
        t <- mod_2096.get(3);
        mod_2097.put(0, t);
    endrule
    rule rule_2728;
        ChannelMessage t;
        t <- mod_2128.get(0);
        mod_2127.put(0, t);
    endrule
    rule rule_2729;
        ChannelMessage t;
        t <- mod_2109.get(0);
        mod_2109.put(1, t);
    endrule
    rule rule_2730;
        ChannelMessage t;
        t <- mod_2131.get(1);
        mod_2095.put(1, t);
    endrule
    rule rule_2731;
        ChannelMessage t;
        t <- mod_2125.get(0);
        mod_2126.put(0, t);
    endrule
    rule rule_2732;
        ChannelMessage t;
        t <- mod_2103.get(1);
        mod_2104.put(0, t);
    endrule
    rule rule_2733;
        ChannelMessage t;
        t <- mod_2113.get(0);
        mod_2111.put(0, t);
    endrule
    rule rule_2734;
        ChannelMessage t;
        t <- mod_2103.get(0);
        mod_2115.put(0, t);
    endrule
    rule rule_2735;
        ChannelMessage t;
        t <- mod_2120.get(0);
        mod_2119.put(1, t);
    endrule
    rule rule_2736;
        ChannelMessage t;
        t <- mod_2094.get(0);
        mod_2095.put(0, t);
    endrule
    rule rule_2737;
        ChannelMessage t;
        t <- mod_2127.get(0);
        mod_2125.put(0, t);
    endrule
    rule rule_2738;
        ChannelMessage t;
        t <- mod_2119.get(0);
        mod_2120.put(0, t);
    endrule
    rule rule_2739;
        ChannelMessage t;
        t <- mod_2123.get(1);
        mod_2118.put(0, t);
    endrule
    rule rule_2740;
        ChannelMessage t;
        t <- mod_2095.get(0);
        mod_2131.put(0, t);
    endrule
    rule rule_2741;
        ChannelMessage t;
        t <- mod_2097.get(0);
        mod_2130.put(0, t);
    endrule
    rule rule_2742;
        ChannelMessage t;
        t <- mod_2110.get(1);
        mod_2106.put(1, t);
    endrule
    rule rule_2743;
        ChannelMessage t;
        t <- mod_2093.get(0);
        mod_2094.put(0, t);
    endrule
    rule rule_2744;
        ChannelMessage t;
        t <- mod_2125.get(1);
        mod_2100.put(1, t);
    endrule
    rule rule_2745;
        ChannelMessage t;
        t <- mod_2100.get(0);
        mod_2101.put(0, t);
    endrule
    rule rule_2746;
        ChannelMessage t;
        t <- mod_2115.get(0);
        mod_2103.put(1, t);
    endrule
    rule rule_2747;
        ChannelMessage t;
        t <- mod_2131.get(0);
        mod_2131.put(1, t);
    endrule
    rule rule_2748;
        ChannelMessage t;
        t <- mod_2095.get(1);
        mod_2096.put(0, t);
    endrule
    rule rule_2749;
        ChannelMessage t;
        t <- mod_2117.get(0);
        mod_2116.put(0, t);
    endrule
    rule rule_2750;
        ChannelMessage t;
        t <- mod_2118.get(0);
        mod_2117.put(0, t);
    endrule
    rule rule_2751;
        ChannelMessage t;
        t <- mod_2107.get(0);
        mod_2109.put(0, t);
    endrule
    rule rule_2752;
        ChannelMessage t;
        t <- mod_2123.get(0);
        mod_2124.put(0, t);
    endrule
    rule rule_2753;
        ChannelMessage t;
        t <- mod_2110.get(0);
        mod_2110.put(1, t);
    endrule
    rule rule_2754;
        ChannelMessage t;
        t <- mod_2105.get(0);
        mod_2106.put(0, t);
    endrule
    rule rule_2755;
        ChannelMessage t;
        t <- mod_2098.get(1);
        mod_2099.put(0, t);
    endrule
    rule rule_2756;
        ChannelMessage t;
        t <- mod_2104.get(0);
        mod_2105.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2092.put(0, t);
        end
        if (i == 1) begin
            mod_2108.put(0, t);
        end
        if (i == 2) begin
            mod_2114.put(0, t);
        end
        if (i == 3) begin
            mod_2122.put(0, t);
        end
        if (i == 4) begin
            mod_2128.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_2096.get(0);
        end
        if (i == 0) begin
            t <- mod_2096.get(1);
        end
        if (i == 1) begin
            t <- mod_2096.get(2);
        end
        if (i == 2) begin
            t <- mod_2108.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6086 (Operation_IFC);
    Operation_IFC mod_2133_inner <- mkReshape(2, 64);
    Operation_IFC mod_2133 <- mkDebugOperation(mod_2133_inner, "mod_2133");
    Operation_IFC mod_2134_inner <- mkFlatten(1);
    Operation_IFC mod_2134 <- mkDebugOperation(mod_2134_inner, "mod_2134");
    Operation_IFC mod_2135_inner <- mkFlatten(2);
    Operation_IFC mod_2135 <- mkDebugOperation(mod_2135_inner, "mod_2135");
    Operation_IFC mod_2136_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2136 <- mkDebugOperation(mod_2136_inner, "mod_2136");
    Broadcast_IFC#(4) mod_2137_inner <- mkBroadcast(4);
    Operation_IFC mod_2137 <- mkDebugOperation(mod_2137_inner.op, "mod_2137");
    PMU_IFC mod_2138_bufferize <- mkPMU(2);
    Operation_IFC mod_2138_inner = mod_2138_bufferize.operation;
    Operation_IFC mod_2138 <- mkDebugOperation(mod_2138_inner, "mod_2138");
    Broadcast_IFC#(2) mod_2139_inner <- mkBroadcast(2);
    Operation_IFC mod_2139 <- mkDebugOperation(mod_2139_inner.op, "mod_2139");
    PMU_IFC mod_2140_bufferize <- mkPMU(1);
    Operation_IFC mod_2140_inner = mod_2140_bufferize.operation;
    Operation_IFC mod_2140 <- mkDebugOperation(mod_2140_inner, "mod_2140");
    Operation_IFC mod_2141_inner <- mkBinaryMap(1104, matmul_t_tile);
    Operation_IFC mod_2141 <- mkDebugOperation(mod_2141_inner, "mod_2141");
    Operation_IFC mod_2142_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2142 <- mkDebugOperation(mod_2142_inner, "mod_2142");
    Operation_IFC mod_2143_inner <- mkBinaryMap(1872, mul_tile);
    Operation_IFC mod_2143 <- mkDebugOperation(mod_2143_inner, "mod_2143");
    PMU_IFC mod_2144_bufferize <- mkPMU(1);
    Operation_IFC mod_2144_inner = mod_2144_bufferize.operation;
    Operation_IFC mod_2144 <- mkDebugOperation(mod_2144_inner, "mod_2144");
    Operation_IFC mod_2145_inner <- mkBinaryMap(2459, matmul_t_tile);
    Operation_IFC mod_2145 <- mkDebugOperation(mod_2145_inner, "mod_2145");
    Operation_IFC mod_2146_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2146 <- mkDebugOperation(mod_2146_inner, "mod_2146");
    Operation_IFC mod_2147_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2147 <- mkDebugOperation(mod_2147_inner, "mod_2147");
    Operation_IFC mod_2148_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2148 <- mkDebugOperation(mod_2148_inner, "mod_2148");
    Operation_IFC mod_2149_inner <- mkBinaryMap(2771, mul_tile);
    Operation_IFC mod_2149 <- mkDebugOperation(mod_2149_inner, "mod_2149");
    PMU_IFC mod_2150_bufferize <- mkPMU(1);
    Operation_IFC mod_2150_inner = mod_2150_bufferize.operation;
    Operation_IFC mod_2150 <- mkDebugOperation(mod_2150_inner, "mod_2150");
    PMU_IFC mod_2151_bufferize <- mkPMU(2);
    Operation_IFC mod_2151_inner = mod_2151_bufferize.operation;
    Operation_IFC mod_2151 <- mkDebugOperation(mod_2151_inner, "mod_2151");
    PMU_IFC mod_2152_bufferize <- mkPMU(2);
    Operation_IFC mod_2152_inner = mod_2152_bufferize.operation;
    Operation_IFC mod_2152 <- mkDebugOperation(mod_2152_inner, "mod_2152");
    Operation_IFC mod_2153_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2153 <- mkDebugOperation(mod_2153_inner, "mod_2153");
    Operation_IFC mod_2154_inner <- mkFlatten(1);
    Operation_IFC mod_2154 <- mkDebugOperation(mod_2154_inner, "mod_2154");
    Operation_IFC mod_2155_inner <- mkFlatten(0);
    Operation_IFC mod_2155 <- mkDebugOperation(mod_2155_inner, "mod_2155");
    Operation_IFC mod_2156_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2156 <- mkDebugOperation(mod_2156_inner, "mod_2156");
    Operation_IFC mod_2157_inner <- mkUnaryMap(1744, silu_tile);
    Operation_IFC mod_2157 <- mkDebugOperation(mod_2157_inner, "mod_2157");
    Operation_IFC mod_2158_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2158 <- mkDebugOperation(mod_2158_inner, "mod_2158");
    Operation_IFC mod_2159_inner <- mkBinaryMap(1616, matmul_t_tile);
    Operation_IFC mod_2159 <- mkDebugOperation(mod_2159_inner, "mod_2159");
    PMU_IFC mod_2160_bufferize <- mkPMU(2);
    Operation_IFC mod_2160_inner = mod_2160_bufferize.operation;
    Operation_IFC mod_2160 <- mkDebugOperation(mod_2160_inner, "mod_2160");
    Operation_IFC mod_2161_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2161 <- mkDebugOperation(mod_2161_inner, "mod_2161");
    Operation_IFC mod_2162_inner <- mkFlatten(1);
    Operation_IFC mod_2162 <- mkDebugOperation(mod_2162_inner, "mod_2162");
    Operation_IFC mod_2163_inner <- mkFlatten(0);
    Operation_IFC mod_2163 <- mkDebugOperation(mod_2163_inner, "mod_2163");
    PMU_IFC mod_2164_bufferize <- mkPMU(1);
    Operation_IFC mod_2164_inner = mod_2164_bufferize.operation;
    Operation_IFC mod_2164 <- mkDebugOperation(mod_2164_inner, "mod_2164");
    Operation_IFC mod_2165_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2165 <- mkDebugOperation(mod_2165_inner, "mod_2165");
    PMU_IFC mod_2166_bufferize <- mkPMU(2);
    Operation_IFC mod_2166_inner = mod_2166_bufferize.operation;
    Operation_IFC mod_2166 <- mkDebugOperation(mod_2166_inner, "mod_2166");
    Operation_IFC mod_2167_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2167 <- mkDebugOperation(mod_2167_inner, "mod_2167");
    Operation_IFC mod_2168_inner <- mkFlatten(1);
    Operation_IFC mod_2168 <- mkDebugOperation(mod_2168_inner, "mod_2168");
    Operation_IFC mod_2169_inner <- mkFlatten(0);
    Operation_IFC mod_2169 <- mkDebugOperation(mod_2169_inner, "mod_2169");
    Operation_IFC mod_2170_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2170 <- mkDebugOperation(mod_2170_inner, "mod_2170");
    Operation_IFC mod_2171_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2171 <- mkDebugOperation(mod_2171_inner, "mod_2171");
    PMU_IFC mod_2172_bufferize <- mkPMU(2);
    Operation_IFC mod_2172_inner = mod_2172_bufferize.operation;
    Operation_IFC mod_2172 <- mkDebugOperation(mod_2172_inner, "mod_2172");
    rule rule_2757;
        ChannelMessage t;
        t <- mod_2166.get(1);
        mod_2141.put(1, t);
    endrule
    rule rule_2758;
        ChannelMessage t;
        t <- mod_2172.get(0);
        mod_2172.put(1, t);
    endrule
    rule rule_2759;
        ChannelMessage t;
        t <- mod_2142.get(0);
        mod_2143.put(0, t);
    endrule
    rule rule_2760;
        ChannelMessage t;
        t <- mod_2169.get(0);
        mod_2168.put(0, t);
    endrule
    rule rule_2761;
        ChannelMessage t;
        t <- mod_2157.get(0);
        mod_2143.put(1, t);
    endrule
    rule rule_2762;
        ChannelMessage t;
        t <- mod_2144.get(1);
        mod_2145.put(0, t);
    endrule
    rule rule_2763;
        ChannelMessage t;
        t <- mod_2160.get(1);
        mod_2159.put(1, t);
    endrule
    rule rule_2764;
        ChannelMessage t;
        t <- mod_2166.get(0);
        mod_2167.put(0, t);
    endrule
    rule rule_2765;
        ChannelMessage t;
        t <- mod_2134.get(0);
        mod_2135.put(0, t);
    endrule
    rule rule_2766;
        ChannelMessage t;
        t <- mod_2165.get(0);
        mod_2164.put(1, t);
    endrule
    rule rule_2767;
        ChannelMessage t;
        t <- mod_2138.get(1);
        mod_2139.put(0, t);
    endrule
    rule rule_2768;
        ChannelMessage t;
        t <- mod_2140.get(0);
        mod_2170.put(0, t);
    endrule
    rule rule_2769;
        ChannelMessage t;
        t <- mod_2144.get(0);
        mod_2156.put(0, t);
    endrule
    rule rule_2770;
        ChannelMessage t;
        t <- mod_2136.get(0);
        mod_2172.put(0, t);
    endrule
    rule rule_2771;
        ChannelMessage t;
        t <- mod_2139.get(1);
        mod_2140.put(0, t);
    endrule
    rule rule_2772;
        ChannelMessage t;
        t <- mod_2156.get(0);
        mod_2144.put(1, t);
    endrule
    rule rule_2773;
        ChannelMessage t;
        t <- mod_2147.get(0);
        mod_2151.put(0, t);
    endrule
    rule rule_2774;
        ChannelMessage t;
        t <- mod_2136.get(1);
        mod_2137.put(0, t);
    endrule
    rule rule_2775;
        ChannelMessage t;
        t <- mod_2158.get(0);
        mod_2157.put(0, t);
    endrule
    rule rule_2776;
        ChannelMessage t;
        t <- mod_2152.get(0);
        mod_2153.put(0, t);
    endrule
    rule rule_2777;
        ChannelMessage t;
        t <- mod_2159.get(0);
        mod_2158.put(0, t);
    endrule
    rule rule_2778;
        ChannelMessage t;
        t <- mod_2170.get(0);
        mod_2140.put(1, t);
    endrule
    rule rule_2779;
        ChannelMessage t;
        t <- mod_2151.get(1);
        mod_2147.put(1, t);
    endrule
    rule rule_2780;
        ChannelMessage t;
        t <- mod_2155.get(0);
        mod_2154.put(0, t);
    endrule
    rule rule_2781;
        ChannelMessage t;
        t <- mod_2163.get(0);
        mod_2162.put(0, t);
    endrule
    rule rule_2782;
        ChannelMessage t;
        t <- mod_2151.get(0);
        mod_2151.put(1, t);
    endrule
    rule rule_2783;
        ChannelMessage t;
        t <- mod_2147.get(1);
        mod_2148.put(0, t);
    endrule
    rule rule_2784;
        ChannelMessage t;
        t <- mod_2133.get(0);
        mod_2134.put(0, t);
    endrule
    rule rule_2785;
        ChannelMessage t;
        t <- mod_2139.get(0);
        mod_2164.put(0, t);
    endrule
    rule rule_2786;
        ChannelMessage t;
        t <- mod_2148.get(0);
        mod_2150.put(0, t);
    endrule
    rule rule_2787;
        ChannelMessage t;
        t <- mod_2140.get(1);
        mod_2141.put(0, t);
    endrule
    rule rule_2788;
        ChannelMessage t;
        t <- mod_2150.get(1);
        mod_2148.put(1, t);
    endrule
    rule rule_2789;
        ChannelMessage t;
        t <- mod_2138.get(0);
        mod_2171.put(0, t);
    endrule
    rule rule_2790;
        ChannelMessage t;
        t <- mod_2172.get(1);
        mod_2136.put(1, t);
    endrule
    rule rule_2791;
        ChannelMessage t;
        t <- mod_2145.get(0);
        mod_2146.put(0, t);
    endrule
    rule rule_2792;
        ChannelMessage t;
        t <- mod_2161.get(0);
        mod_2160.put(1, t);
    endrule
    rule rule_2793;
        ChannelMessage t;
        t <- mod_2164.get(1);
        mod_2159.put(0, t);
    endrule
    rule rule_2794;
        ChannelMessage t;
        t <- mod_2160.get(0);
        mod_2161.put(0, t);
    endrule
    rule rule_2795;
        ChannelMessage t;
        t <- mod_2164.get(0);
        mod_2165.put(0, t);
    endrule
    rule rule_2796;
        ChannelMessage t;
        t <- mod_2135.get(0);
        mod_2136.put(0, t);
    endrule
    rule rule_2797;
        ChannelMessage t;
        t <- mod_2171.get(0);
        mod_2138.put(1, t);
    endrule
    rule rule_2798;
        ChannelMessage t;
        t <- mod_2167.get(0);
        mod_2166.put(1, t);
    endrule
    rule rule_2799;
        ChannelMessage t;
        t <- mod_2143.get(0);
        mod_2144.put(0, t);
    endrule
    rule rule_2800;
        ChannelMessage t;
        t <- mod_2162.get(0);
        mod_2160.put(0, t);
    endrule
    rule rule_2801;
        ChannelMessage t;
        t <- mod_2150.get(0);
        mod_2150.put(1, t);
    endrule
    rule rule_2802;
        ChannelMessage t;
        t <- mod_2153.get(0);
        mod_2152.put(1, t);
    endrule
    rule rule_2803;
        ChannelMessage t;
        t <- mod_2154.get(0);
        mod_2152.put(0, t);
    endrule
    rule rule_2804;
        ChannelMessage t;
        t <- mod_2141.get(0);
        mod_2142.put(0, t);
    endrule
    rule rule_2805;
        ChannelMessage t;
        t <- mod_2152.get(1);
        mod_2145.put(1, t);
    endrule
    rule rule_2806;
        ChannelMessage t;
        t <- mod_2137.get(3);
        mod_2138.put(0, t);
    endrule
    rule rule_2807;
        ChannelMessage t;
        t <- mod_2168.get(0);
        mod_2166.put(0, t);
    endrule
    rule rule_2808;
        ChannelMessage t;
        t <- mod_2146.get(0);
        mod_2147.put(0, t);
    endrule
    rule rule_2809;
        ChannelMessage t;
        t <- mod_2148.get(1);
        mod_2149.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2133.put(0, t);
        end
        if (i == 1) begin
            mod_2149.put(0, t);
        end
        if (i == 2) begin
            mod_2155.put(0, t);
        end
        if (i == 3) begin
            mod_2163.put(0, t);
        end
        if (i == 4) begin
            mod_2169.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_2137.get(0);
        end
        if (i == 3) begin
            t <- mod_2137.get(1);
        end
        if (i == 0) begin
            t <- mod_2137.get(2);
        end
        if (i == 2) begin
            t <- mod_2149.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6087 (Operation_IFC);
    Operation_IFC mod_2174_inner <- mkReshape(2, 64);
    Operation_IFC mod_2174 <- mkDebugOperation(mod_2174_inner, "mod_2174");
    Operation_IFC mod_2175_inner <- mkFlatten(1);
    Operation_IFC mod_2175 <- mkDebugOperation(mod_2175_inner, "mod_2175");
    Operation_IFC mod_2176_inner <- mkFlatten(2);
    Operation_IFC mod_2176 <- mkDebugOperation(mod_2176_inner, "mod_2176");
    Operation_IFC mod_2177_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2177 <- mkDebugOperation(mod_2177_inner, "mod_2177");
    Broadcast_IFC#(4) mod_2178_inner <- mkBroadcast(4);
    Operation_IFC mod_2178 <- mkDebugOperation(mod_2178_inner.op, "mod_2178");
    PMU_IFC mod_2179_bufferize <- mkPMU(2);
    Operation_IFC mod_2179_inner = mod_2179_bufferize.operation;
    Operation_IFC mod_2179 <- mkDebugOperation(mod_2179_inner, "mod_2179");
    Broadcast_IFC#(2) mod_2180_inner <- mkBroadcast(2);
    Operation_IFC mod_2180 <- mkDebugOperation(mod_2180_inner.op, "mod_2180");
    PMU_IFC mod_2181_bufferize <- mkPMU(1);
    Operation_IFC mod_2181_inner = mod_2181_bufferize.operation;
    Operation_IFC mod_2181 <- mkDebugOperation(mod_2181_inner, "mod_2181");
    Operation_IFC mod_2182_inner <- mkBinaryMap(1103, matmul_t_tile);
    Operation_IFC mod_2182 <- mkDebugOperation(mod_2182_inner, "mod_2182");
    Operation_IFC mod_2183_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2183 <- mkDebugOperation(mod_2183_inner, "mod_2183");
    Operation_IFC mod_2184_inner <- mkBinaryMap(1871, mul_tile);
    Operation_IFC mod_2184 <- mkDebugOperation(mod_2184_inner, "mod_2184");
    PMU_IFC mod_2185_bufferize <- mkPMU(1);
    Operation_IFC mod_2185_inner = mod_2185_bufferize.operation;
    Operation_IFC mod_2185 <- mkDebugOperation(mod_2185_inner, "mod_2185");
    Operation_IFC mod_2186_inner <- mkBinaryMap(2457, matmul_t_tile);
    Operation_IFC mod_2186 <- mkDebugOperation(mod_2186_inner, "mod_2186");
    Operation_IFC mod_2187_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2187 <- mkDebugOperation(mod_2187_inner, "mod_2187");
    Operation_IFC mod_2188_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2188 <- mkDebugOperation(mod_2188_inner, "mod_2188");
    Operation_IFC mod_2189_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2189 <- mkDebugOperation(mod_2189_inner, "mod_2189");
    Operation_IFC mod_2190_inner <- mkBinaryMap(2770, mul_tile);
    Operation_IFC mod_2190 <- mkDebugOperation(mod_2190_inner, "mod_2190");
    PMU_IFC mod_2191_bufferize <- mkPMU(1);
    Operation_IFC mod_2191_inner = mod_2191_bufferize.operation;
    Operation_IFC mod_2191 <- mkDebugOperation(mod_2191_inner, "mod_2191");
    PMU_IFC mod_2192_bufferize <- mkPMU(2);
    Operation_IFC mod_2192_inner = mod_2192_bufferize.operation;
    Operation_IFC mod_2192 <- mkDebugOperation(mod_2192_inner, "mod_2192");
    PMU_IFC mod_2193_bufferize <- mkPMU(2);
    Operation_IFC mod_2193_inner = mod_2193_bufferize.operation;
    Operation_IFC mod_2193 <- mkDebugOperation(mod_2193_inner, "mod_2193");
    Operation_IFC mod_2194_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2194 <- mkDebugOperation(mod_2194_inner, "mod_2194");
    Operation_IFC mod_2195_inner <- mkFlatten(1);
    Operation_IFC mod_2195 <- mkDebugOperation(mod_2195_inner, "mod_2195");
    Operation_IFC mod_2196_inner <- mkFlatten(0);
    Operation_IFC mod_2196 <- mkDebugOperation(mod_2196_inner, "mod_2196");
    Operation_IFC mod_2197_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2197 <- mkDebugOperation(mod_2197_inner, "mod_2197");
    Operation_IFC mod_2198_inner <- mkUnaryMap(1743, silu_tile);
    Operation_IFC mod_2198 <- mkDebugOperation(mod_2198_inner, "mod_2198");
    Operation_IFC mod_2199_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2199 <- mkDebugOperation(mod_2199_inner, "mod_2199");
    Operation_IFC mod_2200_inner <- mkBinaryMap(1615, matmul_t_tile);
    Operation_IFC mod_2200 <- mkDebugOperation(mod_2200_inner, "mod_2200");
    PMU_IFC mod_2201_bufferize <- mkPMU(2);
    Operation_IFC mod_2201_inner = mod_2201_bufferize.operation;
    Operation_IFC mod_2201 <- mkDebugOperation(mod_2201_inner, "mod_2201");
    Operation_IFC mod_2202_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2202 <- mkDebugOperation(mod_2202_inner, "mod_2202");
    Operation_IFC mod_2203_inner <- mkFlatten(1);
    Operation_IFC mod_2203 <- mkDebugOperation(mod_2203_inner, "mod_2203");
    Operation_IFC mod_2204_inner <- mkFlatten(0);
    Operation_IFC mod_2204 <- mkDebugOperation(mod_2204_inner, "mod_2204");
    PMU_IFC mod_2205_bufferize <- mkPMU(1);
    Operation_IFC mod_2205_inner = mod_2205_bufferize.operation;
    Operation_IFC mod_2205 <- mkDebugOperation(mod_2205_inner, "mod_2205");
    Operation_IFC mod_2206_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2206 <- mkDebugOperation(mod_2206_inner, "mod_2206");
    PMU_IFC mod_2207_bufferize <- mkPMU(2);
    Operation_IFC mod_2207_inner = mod_2207_bufferize.operation;
    Operation_IFC mod_2207 <- mkDebugOperation(mod_2207_inner, "mod_2207");
    Operation_IFC mod_2208_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2208 <- mkDebugOperation(mod_2208_inner, "mod_2208");
    Operation_IFC mod_2209_inner <- mkFlatten(1);
    Operation_IFC mod_2209 <- mkDebugOperation(mod_2209_inner, "mod_2209");
    Operation_IFC mod_2210_inner <- mkFlatten(0);
    Operation_IFC mod_2210 <- mkDebugOperation(mod_2210_inner, "mod_2210");
    Operation_IFC mod_2211_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2211 <- mkDebugOperation(mod_2211_inner, "mod_2211");
    Operation_IFC mod_2212_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2212 <- mkDebugOperation(mod_2212_inner, "mod_2212");
    PMU_IFC mod_2213_bufferize <- mkPMU(2);
    Operation_IFC mod_2213_inner = mod_2213_bufferize.operation;
    Operation_IFC mod_2213 <- mkDebugOperation(mod_2213_inner, "mod_2213");
    rule rule_2810;
        ChannelMessage t;
        t <- mod_2213.get(1);
        mod_2177.put(1, t);
    endrule
    rule rule_2811;
        ChannelMessage t;
        t <- mod_2210.get(0);
        mod_2209.put(0, t);
    endrule
    rule rule_2812;
        ChannelMessage t;
        t <- mod_2188.get(1);
        mod_2189.put(0, t);
    endrule
    rule rule_2813;
        ChannelMessage t;
        t <- mod_2203.get(0);
        mod_2201.put(0, t);
    endrule
    rule rule_2814;
        ChannelMessage t;
        t <- mod_2186.get(0);
        mod_2187.put(0, t);
    endrule
    rule rule_2815;
        ChannelMessage t;
        t <- mod_2213.get(0);
        mod_2213.put(1, t);
    endrule
    rule rule_2816;
        ChannelMessage t;
        t <- mod_2192.get(1);
        mod_2188.put(1, t);
    endrule
    rule rule_2817;
        ChannelMessage t;
        t <- mod_2183.get(0);
        mod_2184.put(0, t);
    endrule
    rule rule_2818;
        ChannelMessage t;
        t <- mod_2207.get(0);
        mod_2208.put(0, t);
    endrule
    rule rule_2819;
        ChannelMessage t;
        t <- mod_2208.get(0);
        mod_2207.put(1, t);
    endrule
    rule rule_2820;
        ChannelMessage t;
        t <- mod_2199.get(0);
        mod_2198.put(0, t);
    endrule
    rule rule_2821;
        ChannelMessage t;
        t <- mod_2198.get(0);
        mod_2184.put(1, t);
    endrule
    rule rule_2822;
        ChannelMessage t;
        t <- mod_2181.get(1);
        mod_2182.put(0, t);
    endrule
    rule rule_2823;
        ChannelMessage t;
        t <- mod_2201.get(1);
        mod_2200.put(1, t);
    endrule
    rule rule_2824;
        ChannelMessage t;
        t <- mod_2192.get(0);
        mod_2192.put(1, t);
    endrule
    rule rule_2825;
        ChannelMessage t;
        t <- mod_2200.get(0);
        mod_2199.put(0, t);
    endrule
    rule rule_2826;
        ChannelMessage t;
        t <- mod_2189.get(1);
        mod_2190.put(1, t);
    endrule
    rule rule_2827;
        ChannelMessage t;
        t <- mod_2189.get(0);
        mod_2191.put(0, t);
    endrule
    rule rule_2828;
        ChannelMessage t;
        t <- mod_2205.get(0);
        mod_2206.put(0, t);
    endrule
    rule rule_2829;
        ChannelMessage t;
        t <- mod_2193.get(1);
        mod_2186.put(1, t);
    endrule
    rule rule_2830;
        ChannelMessage t;
        t <- mod_2207.get(1);
        mod_2182.put(1, t);
    endrule
    rule rule_2831;
        ChannelMessage t;
        t <- mod_2194.get(0);
        mod_2193.put(1, t);
    endrule
    rule rule_2832;
        ChannelMessage t;
        t <- mod_2204.get(0);
        mod_2203.put(0, t);
    endrule
    rule rule_2833;
        ChannelMessage t;
        t <- mod_2177.get(0);
        mod_2213.put(0, t);
    endrule
    rule rule_2834;
        ChannelMessage t;
        t <- mod_2174.get(0);
        mod_2175.put(0, t);
    endrule
    rule rule_2835;
        ChannelMessage t;
        t <- mod_2179.get(1);
        mod_2180.put(0, t);
    endrule
    rule rule_2836;
        ChannelMessage t;
        t <- mod_2195.get(0);
        mod_2193.put(0, t);
    endrule
    rule rule_2837;
        ChannelMessage t;
        t <- mod_2191.get(1);
        mod_2189.put(1, t);
    endrule
    rule rule_2838;
        ChannelMessage t;
        t <- mod_2209.get(0);
        mod_2207.put(0, t);
    endrule
    rule rule_2839;
        ChannelMessage t;
        t <- mod_2176.get(0);
        mod_2177.put(0, t);
    endrule
    rule rule_2840;
        ChannelMessage t;
        t <- mod_2177.get(1);
        mod_2178.put(0, t);
    endrule
    rule rule_2841;
        ChannelMessage t;
        t <- mod_2206.get(0);
        mod_2205.put(1, t);
    endrule
    rule rule_2842;
        ChannelMessage t;
        t <- mod_2202.get(0);
        mod_2201.put(1, t);
    endrule
    rule rule_2843;
        ChannelMessage t;
        t <- mod_2212.get(0);
        mod_2179.put(1, t);
    endrule
    rule rule_2844;
        ChannelMessage t;
        t <- mod_2180.get(0);
        mod_2205.put(0, t);
    endrule
    rule rule_2845;
        ChannelMessage t;
        t <- mod_2196.get(0);
        mod_2195.put(0, t);
    endrule
    rule rule_2846;
        ChannelMessage t;
        t <- mod_2175.get(0);
        mod_2176.put(0, t);
    endrule
    rule rule_2847;
        ChannelMessage t;
        t <- mod_2197.get(0);
        mod_2185.put(1, t);
    endrule
    rule rule_2848;
        ChannelMessage t;
        t <- mod_2178.get(3);
        mod_2179.put(0, t);
    endrule
    rule rule_2849;
        ChannelMessage t;
        t <- mod_2182.get(0);
        mod_2183.put(0, t);
    endrule
    rule rule_2850;
        ChannelMessage t;
        t <- mod_2184.get(0);
        mod_2185.put(0, t);
    endrule
    rule rule_2851;
        ChannelMessage t;
        t <- mod_2185.get(0);
        mod_2197.put(0, t);
    endrule
    rule rule_2852;
        ChannelMessage t;
        t <- mod_2205.get(1);
        mod_2200.put(0, t);
    endrule
    rule rule_2853;
        ChannelMessage t;
        t <- mod_2211.get(0);
        mod_2181.put(1, t);
    endrule
    rule rule_2854;
        ChannelMessage t;
        t <- mod_2180.get(1);
        mod_2181.put(0, t);
    endrule
    rule rule_2855;
        ChannelMessage t;
        t <- mod_2193.get(0);
        mod_2194.put(0, t);
    endrule
    rule rule_2856;
        ChannelMessage t;
        t <- mod_2181.get(0);
        mod_2211.put(0, t);
    endrule
    rule rule_2857;
        ChannelMessage t;
        t <- mod_2185.get(1);
        mod_2186.put(0, t);
    endrule
    rule rule_2858;
        ChannelMessage t;
        t <- mod_2191.get(0);
        mod_2191.put(1, t);
    endrule
    rule rule_2859;
        ChannelMessage t;
        t <- mod_2179.get(0);
        mod_2212.put(0, t);
    endrule
    rule rule_2860;
        ChannelMessage t;
        t <- mod_2187.get(0);
        mod_2188.put(0, t);
    endrule
    rule rule_2861;
        ChannelMessage t;
        t <- mod_2188.get(0);
        mod_2192.put(0, t);
    endrule
    rule rule_2862;
        ChannelMessage t;
        t <- mod_2201.get(0);
        mod_2202.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2174.put(0, t);
        end
        if (i == 1) begin
            mod_2190.put(0, t);
        end
        if (i == 2) begin
            mod_2196.put(0, t);
        end
        if (i == 3) begin
            mod_2204.put(0, t);
        end
        if (i == 4) begin
            mod_2210.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_2178.get(0);
        end
        if (i == 3) begin
            t <- mod_2178.get(1);
        end
        if (i == 0) begin
            t <- mod_2178.get(2);
        end
        if (i == 2) begin
            t <- mod_2190.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6088 (Operation_IFC);
    Operation_IFC mod_2215_inner <- mkReshape(2, 64);
    Operation_IFC mod_2215 <- mkDebugOperation(mod_2215_inner, "mod_2215");
    Operation_IFC mod_2216_inner <- mkFlatten(1);
    Operation_IFC mod_2216 <- mkDebugOperation(mod_2216_inner, "mod_2216");
    Operation_IFC mod_2217_inner <- mkFlatten(2);
    Operation_IFC mod_2217 <- mkDebugOperation(mod_2217_inner, "mod_2217");
    Operation_IFC mod_2218_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2218 <- mkDebugOperation(mod_2218_inner, "mod_2218");
    Broadcast_IFC#(4) mod_2219_inner <- mkBroadcast(4);
    Operation_IFC mod_2219 <- mkDebugOperation(mod_2219_inner.op, "mod_2219");
    PMU_IFC mod_2220_bufferize <- mkPMU(2);
    Operation_IFC mod_2220_inner = mod_2220_bufferize.operation;
    Operation_IFC mod_2220 <- mkDebugOperation(mod_2220_inner, "mod_2220");
    Broadcast_IFC#(2) mod_2221_inner <- mkBroadcast(2);
    Operation_IFC mod_2221 <- mkDebugOperation(mod_2221_inner.op, "mod_2221");
    PMU_IFC mod_2222_bufferize <- mkPMU(1);
    Operation_IFC mod_2222_inner = mod_2222_bufferize.operation;
    Operation_IFC mod_2222 <- mkDebugOperation(mod_2222_inner, "mod_2222");
    Operation_IFC mod_2223_inner <- mkBinaryMap(1102, matmul_t_tile);
    Operation_IFC mod_2223 <- mkDebugOperation(mod_2223_inner, "mod_2223");
    Operation_IFC mod_2224_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2224 <- mkDebugOperation(mod_2224_inner, "mod_2224");
    Operation_IFC mod_2225_inner <- mkBinaryMap(1870, mul_tile);
    Operation_IFC mod_2225 <- mkDebugOperation(mod_2225_inner, "mod_2225");
    PMU_IFC mod_2226_bufferize <- mkPMU(1);
    Operation_IFC mod_2226_inner = mod_2226_bufferize.operation;
    Operation_IFC mod_2226 <- mkDebugOperation(mod_2226_inner, "mod_2226");
    Operation_IFC mod_2227_inner <- mkBinaryMap(2455, matmul_t_tile);
    Operation_IFC mod_2227 <- mkDebugOperation(mod_2227_inner, "mod_2227");
    Operation_IFC mod_2228_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2228 <- mkDebugOperation(mod_2228_inner, "mod_2228");
    Operation_IFC mod_2229_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2229 <- mkDebugOperation(mod_2229_inner, "mod_2229");
    Operation_IFC mod_2230_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2230 <- mkDebugOperation(mod_2230_inner, "mod_2230");
    Operation_IFC mod_2231_inner <- mkBinaryMap(2769, mul_tile);
    Operation_IFC mod_2231 <- mkDebugOperation(mod_2231_inner, "mod_2231");
    PMU_IFC mod_2232_bufferize <- mkPMU(1);
    Operation_IFC mod_2232_inner = mod_2232_bufferize.operation;
    Operation_IFC mod_2232 <- mkDebugOperation(mod_2232_inner, "mod_2232");
    PMU_IFC mod_2233_bufferize <- mkPMU(2);
    Operation_IFC mod_2233_inner = mod_2233_bufferize.operation;
    Operation_IFC mod_2233 <- mkDebugOperation(mod_2233_inner, "mod_2233");
    PMU_IFC mod_2234_bufferize <- mkPMU(2);
    Operation_IFC mod_2234_inner = mod_2234_bufferize.operation;
    Operation_IFC mod_2234 <- mkDebugOperation(mod_2234_inner, "mod_2234");
    Operation_IFC mod_2235_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2235 <- mkDebugOperation(mod_2235_inner, "mod_2235");
    Operation_IFC mod_2236_inner <- mkFlatten(1);
    Operation_IFC mod_2236 <- mkDebugOperation(mod_2236_inner, "mod_2236");
    Operation_IFC mod_2237_inner <- mkFlatten(0);
    Operation_IFC mod_2237 <- mkDebugOperation(mod_2237_inner, "mod_2237");
    Operation_IFC mod_2238_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2238 <- mkDebugOperation(mod_2238_inner, "mod_2238");
    Operation_IFC mod_2239_inner <- mkUnaryMap(1742, silu_tile);
    Operation_IFC mod_2239 <- mkDebugOperation(mod_2239_inner, "mod_2239");
    Operation_IFC mod_2240_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2240 <- mkDebugOperation(mod_2240_inner, "mod_2240");
    Operation_IFC mod_2241_inner <- mkBinaryMap(1614, matmul_t_tile);
    Operation_IFC mod_2241 <- mkDebugOperation(mod_2241_inner, "mod_2241");
    PMU_IFC mod_2242_bufferize <- mkPMU(2);
    Operation_IFC mod_2242_inner = mod_2242_bufferize.operation;
    Operation_IFC mod_2242 <- mkDebugOperation(mod_2242_inner, "mod_2242");
    Operation_IFC mod_2243_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2243 <- mkDebugOperation(mod_2243_inner, "mod_2243");
    Operation_IFC mod_2244_inner <- mkFlatten(1);
    Operation_IFC mod_2244 <- mkDebugOperation(mod_2244_inner, "mod_2244");
    Operation_IFC mod_2245_inner <- mkFlatten(0);
    Operation_IFC mod_2245 <- mkDebugOperation(mod_2245_inner, "mod_2245");
    PMU_IFC mod_2246_bufferize <- mkPMU(1);
    Operation_IFC mod_2246_inner = mod_2246_bufferize.operation;
    Operation_IFC mod_2246 <- mkDebugOperation(mod_2246_inner, "mod_2246");
    Operation_IFC mod_2247_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2247 <- mkDebugOperation(mod_2247_inner, "mod_2247");
    PMU_IFC mod_2248_bufferize <- mkPMU(2);
    Operation_IFC mod_2248_inner = mod_2248_bufferize.operation;
    Operation_IFC mod_2248 <- mkDebugOperation(mod_2248_inner, "mod_2248");
    Operation_IFC mod_2249_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2249 <- mkDebugOperation(mod_2249_inner, "mod_2249");
    Operation_IFC mod_2250_inner <- mkFlatten(1);
    Operation_IFC mod_2250 <- mkDebugOperation(mod_2250_inner, "mod_2250");
    Operation_IFC mod_2251_inner <- mkFlatten(0);
    Operation_IFC mod_2251 <- mkDebugOperation(mod_2251_inner, "mod_2251");
    Operation_IFC mod_2252_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2252 <- mkDebugOperation(mod_2252_inner, "mod_2252");
    Operation_IFC mod_2253_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2253 <- mkDebugOperation(mod_2253_inner, "mod_2253");
    PMU_IFC mod_2254_bufferize <- mkPMU(2);
    Operation_IFC mod_2254_inner = mod_2254_bufferize.operation;
    Operation_IFC mod_2254 <- mkDebugOperation(mod_2254_inner, "mod_2254");
    rule rule_2863;
        ChannelMessage t;
        t <- mod_2230.get(1);
        mod_2231.put(1, t);
    endrule
    rule rule_2864;
        ChannelMessage t;
        t <- mod_2218.get(1);
        mod_2219.put(0, t);
    endrule
    rule rule_2865;
        ChannelMessage t;
        t <- mod_2227.get(0);
        mod_2228.put(0, t);
    endrule
    rule rule_2866;
        ChannelMessage t;
        t <- mod_2249.get(0);
        mod_2248.put(1, t);
    endrule
    rule rule_2867;
        ChannelMessage t;
        t <- mod_2225.get(0);
        mod_2226.put(0, t);
    endrule
    rule rule_2868;
        ChannelMessage t;
        t <- mod_2243.get(0);
        mod_2242.put(1, t);
    endrule
    rule rule_2869;
        ChannelMessage t;
        t <- mod_2222.get(1);
        mod_2223.put(0, t);
    endrule
    rule rule_2870;
        ChannelMessage t;
        t <- mod_2215.get(0);
        mod_2216.put(0, t);
    endrule
    rule rule_2871;
        ChannelMessage t;
        t <- mod_2233.get(1);
        mod_2229.put(1, t);
    endrule
    rule rule_2872;
        ChannelMessage t;
        t <- mod_2237.get(0);
        mod_2236.put(0, t);
    endrule
    rule rule_2873;
        ChannelMessage t;
        t <- mod_2220.get(1);
        mod_2221.put(0, t);
    endrule
    rule rule_2874;
        ChannelMessage t;
        t <- mod_2220.get(0);
        mod_2253.put(0, t);
    endrule
    rule rule_2875;
        ChannelMessage t;
        t <- mod_2239.get(0);
        mod_2225.put(1, t);
    endrule
    rule rule_2876;
        ChannelMessage t;
        t <- mod_2221.get(0);
        mod_2246.put(0, t);
    endrule
    rule rule_2877;
        ChannelMessage t;
        t <- mod_2235.get(0);
        mod_2234.put(1, t);
    endrule
    rule rule_2878;
        ChannelMessage t;
        t <- mod_2240.get(0);
        mod_2239.put(0, t);
    endrule
    rule rule_2879;
        ChannelMessage t;
        t <- mod_2254.get(0);
        mod_2254.put(1, t);
    endrule
    rule rule_2880;
        ChannelMessage t;
        t <- mod_2234.get(1);
        mod_2227.put(1, t);
    endrule
    rule rule_2881;
        ChannelMessage t;
        t <- mod_2246.get(0);
        mod_2247.put(0, t);
    endrule
    rule rule_2882;
        ChannelMessage t;
        t <- mod_2219.get(3);
        mod_2220.put(0, t);
    endrule
    rule rule_2883;
        ChannelMessage t;
        t <- mod_2251.get(0);
        mod_2250.put(0, t);
    endrule
    rule rule_2884;
        ChannelMessage t;
        t <- mod_2217.get(0);
        mod_2218.put(0, t);
    endrule
    rule rule_2885;
        ChannelMessage t;
        t <- mod_2234.get(0);
        mod_2235.put(0, t);
    endrule
    rule rule_2886;
        ChannelMessage t;
        t <- mod_2224.get(0);
        mod_2225.put(0, t);
    endrule
    rule rule_2887;
        ChannelMessage t;
        t <- mod_2253.get(0);
        mod_2220.put(1, t);
    endrule
    rule rule_2888;
        ChannelMessage t;
        t <- mod_2254.get(1);
        mod_2218.put(1, t);
    endrule
    rule rule_2889;
        ChannelMessage t;
        t <- mod_2246.get(1);
        mod_2241.put(0, t);
    endrule
    rule rule_2890;
        ChannelMessage t;
        t <- mod_2221.get(1);
        mod_2222.put(0, t);
    endrule
    rule rule_2891;
        ChannelMessage t;
        t <- mod_2229.get(1);
        mod_2230.put(0, t);
    endrule
    rule rule_2892;
        ChannelMessage t;
        t <- mod_2230.get(0);
        mod_2232.put(0, t);
    endrule
    rule rule_2893;
        ChannelMessage t;
        t <- mod_2236.get(0);
        mod_2234.put(0, t);
    endrule
    rule rule_2894;
        ChannelMessage t;
        t <- mod_2223.get(0);
        mod_2224.put(0, t);
    endrule
    rule rule_2895;
        ChannelMessage t;
        t <- mod_2233.get(0);
        mod_2233.put(1, t);
    endrule
    rule rule_2896;
        ChannelMessage t;
        t <- mod_2228.get(0);
        mod_2229.put(0, t);
    endrule
    rule rule_2897;
        ChannelMessage t;
        t <- mod_2244.get(0);
        mod_2242.put(0, t);
    endrule
    rule rule_2898;
        ChannelMessage t;
        t <- mod_2250.get(0);
        mod_2248.put(0, t);
    endrule
    rule rule_2899;
        ChannelMessage t;
        t <- mod_2226.get(0);
        mod_2238.put(0, t);
    endrule
    rule rule_2900;
        ChannelMessage t;
        t <- mod_2216.get(0);
        mod_2217.put(0, t);
    endrule
    rule rule_2901;
        ChannelMessage t;
        t <- mod_2241.get(0);
        mod_2240.put(0, t);
    endrule
    rule rule_2902;
        ChannelMessage t;
        t <- mod_2222.get(0);
        mod_2252.put(0, t);
    endrule
    rule rule_2903;
        ChannelMessage t;
        t <- mod_2242.get(0);
        mod_2243.put(0, t);
    endrule
    rule rule_2904;
        ChannelMessage t;
        t <- mod_2252.get(0);
        mod_2222.put(1, t);
    endrule
    rule rule_2905;
        ChannelMessage t;
        t <- mod_2245.get(0);
        mod_2244.put(0, t);
    endrule
    rule rule_2906;
        ChannelMessage t;
        t <- mod_2226.get(1);
        mod_2227.put(0, t);
    endrule
    rule rule_2907;
        ChannelMessage t;
        t <- mod_2242.get(1);
        mod_2241.put(1, t);
    endrule
    rule rule_2908;
        ChannelMessage t;
        t <- mod_2232.get(1);
        mod_2230.put(1, t);
    endrule
    rule rule_2909;
        ChannelMessage t;
        t <- mod_2248.get(0);
        mod_2249.put(0, t);
    endrule
    rule rule_2910;
        ChannelMessage t;
        t <- mod_2248.get(1);
        mod_2223.put(1, t);
    endrule
    rule rule_2911;
        ChannelMessage t;
        t <- mod_2238.get(0);
        mod_2226.put(1, t);
    endrule
    rule rule_2912;
        ChannelMessage t;
        t <- mod_2229.get(0);
        mod_2233.put(0, t);
    endrule
    rule rule_2913;
        ChannelMessage t;
        t <- mod_2232.get(0);
        mod_2232.put(1, t);
    endrule
    rule rule_2914;
        ChannelMessage t;
        t <- mod_2218.get(0);
        mod_2254.put(0, t);
    endrule
    rule rule_2915;
        ChannelMessage t;
        t <- mod_2247.get(0);
        mod_2246.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2215.put(0, t);
        end
        if (i == 1) begin
            mod_2231.put(0, t);
        end
        if (i == 2) begin
            mod_2237.put(0, t);
        end
        if (i == 3) begin
            mod_2245.put(0, t);
        end
        if (i == 4) begin
            mod_2251.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 2) begin
            t <- mod_2219.get(0);
        end
        if (i == 3) begin
            t <- mod_2219.get(1);
        end
        if (i == 1) begin
            t <- mod_2219.get(2);
        end
        if (i == 0) begin
            t <- mod_2231.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6089 (Operation_IFC);
    Operation_IFC mod_2256_inner <- mkReshape(2, 64);
    Operation_IFC mod_2256 <- mkDebugOperation(mod_2256_inner, "mod_2256");
    Operation_IFC mod_2257_inner <- mkFlatten(1);
    Operation_IFC mod_2257 <- mkDebugOperation(mod_2257_inner, "mod_2257");
    Operation_IFC mod_2258_inner <- mkFlatten(2);
    Operation_IFC mod_2258 <- mkDebugOperation(mod_2258_inner, "mod_2258");
    Operation_IFC mod_2259_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2259 <- mkDebugOperation(mod_2259_inner, "mod_2259");
    Broadcast_IFC#(4) mod_2260_inner <- mkBroadcast(4);
    Operation_IFC mod_2260 <- mkDebugOperation(mod_2260_inner.op, "mod_2260");
    PMU_IFC mod_2261_bufferize <- mkPMU(2);
    Operation_IFC mod_2261_inner = mod_2261_bufferize.operation;
    Operation_IFC mod_2261 <- mkDebugOperation(mod_2261_inner, "mod_2261");
    Broadcast_IFC#(2) mod_2262_inner <- mkBroadcast(2);
    Operation_IFC mod_2262 <- mkDebugOperation(mod_2262_inner.op, "mod_2262");
    PMU_IFC mod_2263_bufferize <- mkPMU(1);
    Operation_IFC mod_2263_inner = mod_2263_bufferize.operation;
    Operation_IFC mod_2263 <- mkDebugOperation(mod_2263_inner, "mod_2263");
    Operation_IFC mod_2264_inner <- mkBinaryMap(1101, matmul_t_tile);
    Operation_IFC mod_2264 <- mkDebugOperation(mod_2264_inner, "mod_2264");
    Operation_IFC mod_2265_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2265 <- mkDebugOperation(mod_2265_inner, "mod_2265");
    Operation_IFC mod_2266_inner <- mkBinaryMap(1869, mul_tile);
    Operation_IFC mod_2266 <- mkDebugOperation(mod_2266_inner, "mod_2266");
    PMU_IFC mod_2267_bufferize <- mkPMU(1);
    Operation_IFC mod_2267_inner = mod_2267_bufferize.operation;
    Operation_IFC mod_2267 <- mkDebugOperation(mod_2267_inner, "mod_2267");
    Operation_IFC mod_2268_inner <- mkBinaryMap(2453, matmul_t_tile);
    Operation_IFC mod_2268 <- mkDebugOperation(mod_2268_inner, "mod_2268");
    Operation_IFC mod_2269_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2269 <- mkDebugOperation(mod_2269_inner, "mod_2269");
    Operation_IFC mod_2270_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2270 <- mkDebugOperation(mod_2270_inner, "mod_2270");
    Operation_IFC mod_2271_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2271 <- mkDebugOperation(mod_2271_inner, "mod_2271");
    Operation_IFC mod_2272_inner <- mkBinaryMap(2768, mul_tile);
    Operation_IFC mod_2272 <- mkDebugOperation(mod_2272_inner, "mod_2272");
    PMU_IFC mod_2273_bufferize <- mkPMU(1);
    Operation_IFC mod_2273_inner = mod_2273_bufferize.operation;
    Operation_IFC mod_2273 <- mkDebugOperation(mod_2273_inner, "mod_2273");
    PMU_IFC mod_2274_bufferize <- mkPMU(2);
    Operation_IFC mod_2274_inner = mod_2274_bufferize.operation;
    Operation_IFC mod_2274 <- mkDebugOperation(mod_2274_inner, "mod_2274");
    PMU_IFC mod_2275_bufferize <- mkPMU(2);
    Operation_IFC mod_2275_inner = mod_2275_bufferize.operation;
    Operation_IFC mod_2275 <- mkDebugOperation(mod_2275_inner, "mod_2275");
    Operation_IFC mod_2276_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2276 <- mkDebugOperation(mod_2276_inner, "mod_2276");
    Operation_IFC mod_2277_inner <- mkFlatten(1);
    Operation_IFC mod_2277 <- mkDebugOperation(mod_2277_inner, "mod_2277");
    Operation_IFC mod_2278_inner <- mkFlatten(0);
    Operation_IFC mod_2278 <- mkDebugOperation(mod_2278_inner, "mod_2278");
    Operation_IFC mod_2279_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2279 <- mkDebugOperation(mod_2279_inner, "mod_2279");
    Operation_IFC mod_2280_inner <- mkUnaryMap(1741, silu_tile);
    Operation_IFC mod_2280 <- mkDebugOperation(mod_2280_inner, "mod_2280");
    Operation_IFC mod_2281_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2281 <- mkDebugOperation(mod_2281_inner, "mod_2281");
    Operation_IFC mod_2282_inner <- mkBinaryMap(1613, matmul_t_tile);
    Operation_IFC mod_2282 <- mkDebugOperation(mod_2282_inner, "mod_2282");
    PMU_IFC mod_2283_bufferize <- mkPMU(2);
    Operation_IFC mod_2283_inner = mod_2283_bufferize.operation;
    Operation_IFC mod_2283 <- mkDebugOperation(mod_2283_inner, "mod_2283");
    Operation_IFC mod_2284_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2284 <- mkDebugOperation(mod_2284_inner, "mod_2284");
    Operation_IFC mod_2285_inner <- mkFlatten(1);
    Operation_IFC mod_2285 <- mkDebugOperation(mod_2285_inner, "mod_2285");
    Operation_IFC mod_2286_inner <- mkFlatten(0);
    Operation_IFC mod_2286 <- mkDebugOperation(mod_2286_inner, "mod_2286");
    PMU_IFC mod_2287_bufferize <- mkPMU(1);
    Operation_IFC mod_2287_inner = mod_2287_bufferize.operation;
    Operation_IFC mod_2287 <- mkDebugOperation(mod_2287_inner, "mod_2287");
    Operation_IFC mod_2288_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2288 <- mkDebugOperation(mod_2288_inner, "mod_2288");
    PMU_IFC mod_2289_bufferize <- mkPMU(2);
    Operation_IFC mod_2289_inner = mod_2289_bufferize.operation;
    Operation_IFC mod_2289 <- mkDebugOperation(mod_2289_inner, "mod_2289");
    Operation_IFC mod_2290_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2290 <- mkDebugOperation(mod_2290_inner, "mod_2290");
    Operation_IFC mod_2291_inner <- mkFlatten(1);
    Operation_IFC mod_2291 <- mkDebugOperation(mod_2291_inner, "mod_2291");
    Operation_IFC mod_2292_inner <- mkFlatten(0);
    Operation_IFC mod_2292 <- mkDebugOperation(mod_2292_inner, "mod_2292");
    Operation_IFC mod_2293_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2293 <- mkDebugOperation(mod_2293_inner, "mod_2293");
    Operation_IFC mod_2294_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2294 <- mkDebugOperation(mod_2294_inner, "mod_2294");
    PMU_IFC mod_2295_bufferize <- mkPMU(2);
    Operation_IFC mod_2295_inner = mod_2295_bufferize.operation;
    Operation_IFC mod_2295 <- mkDebugOperation(mod_2295_inner, "mod_2295");
    rule rule_2916;
        ChannelMessage t;
        t <- mod_2294.get(0);
        mod_2261.put(1, t);
    endrule
    rule rule_2917;
        ChannelMessage t;
        t <- mod_2264.get(0);
        mod_2265.put(0, t);
    endrule
    rule rule_2918;
        ChannelMessage t;
        t <- mod_2287.get(0);
        mod_2288.put(0, t);
    endrule
    rule rule_2919;
        ChannelMessage t;
        t <- mod_2295.get(1);
        mod_2259.put(1, t);
    endrule
    rule rule_2920;
        ChannelMessage t;
        t <- mod_2276.get(0);
        mod_2275.put(1, t);
    endrule
    rule rule_2921;
        ChannelMessage t;
        t <- mod_2283.get(0);
        mod_2284.put(0, t);
    endrule
    rule rule_2922;
        ChannelMessage t;
        t <- mod_2266.get(0);
        mod_2267.put(0, t);
    endrule
    rule rule_2923;
        ChannelMessage t;
        t <- mod_2283.get(1);
        mod_2282.put(1, t);
    endrule
    rule rule_2924;
        ChannelMessage t;
        t <- mod_2263.get(0);
        mod_2293.put(0, t);
    endrule
    rule rule_2925;
        ChannelMessage t;
        t <- mod_2259.get(1);
        mod_2260.put(0, t);
    endrule
    rule rule_2926;
        ChannelMessage t;
        t <- mod_2280.get(0);
        mod_2266.put(1, t);
    endrule
    rule rule_2927;
        ChannelMessage t;
        t <- mod_2278.get(0);
        mod_2277.put(0, t);
    endrule
    rule rule_2928;
        ChannelMessage t;
        t <- mod_2287.get(1);
        mod_2282.put(0, t);
    endrule
    rule rule_2929;
        ChannelMessage t;
        t <- mod_2274.get(0);
        mod_2274.put(1, t);
    endrule
    rule rule_2930;
        ChannelMessage t;
        t <- mod_2256.get(0);
        mod_2257.put(0, t);
    endrule
    rule rule_2931;
        ChannelMessage t;
        t <- mod_2269.get(0);
        mod_2270.put(0, t);
    endrule
    rule rule_2932;
        ChannelMessage t;
        t <- mod_2293.get(0);
        mod_2263.put(1, t);
    endrule
    rule rule_2933;
        ChannelMessage t;
        t <- mod_2295.get(0);
        mod_2295.put(1, t);
    endrule
    rule rule_2934;
        ChannelMessage t;
        t <- mod_2257.get(0);
        mod_2258.put(0, t);
    endrule
    rule rule_2935;
        ChannelMessage t;
        t <- mod_2289.get(1);
        mod_2264.put(1, t);
    endrule
    rule rule_2936;
        ChannelMessage t;
        t <- mod_2292.get(0);
        mod_2291.put(0, t);
    endrule
    rule rule_2937;
        ChannelMessage t;
        t <- mod_2270.get(1);
        mod_2271.put(0, t);
    endrule
    rule rule_2938;
        ChannelMessage t;
        t <- mod_2273.get(1);
        mod_2271.put(1, t);
    endrule
    rule rule_2939;
        ChannelMessage t;
        t <- mod_2270.get(0);
        mod_2274.put(0, t);
    endrule
    rule rule_2940;
        ChannelMessage t;
        t <- mod_2262.get(0);
        mod_2287.put(0, t);
    endrule
    rule rule_2941;
        ChannelMessage t;
        t <- mod_2268.get(0);
        mod_2269.put(0, t);
    endrule
    rule rule_2942;
        ChannelMessage t;
        t <- mod_2286.get(0);
        mod_2285.put(0, t);
    endrule
    rule rule_2943;
        ChannelMessage t;
        t <- mod_2290.get(0);
        mod_2289.put(1, t);
    endrule
    rule rule_2944;
        ChannelMessage t;
        t <- mod_2291.get(0);
        mod_2289.put(0, t);
    endrule
    rule rule_2945;
        ChannelMessage t;
        t <- mod_2259.get(0);
        mod_2295.put(0, t);
    endrule
    rule rule_2946;
        ChannelMessage t;
        t <- mod_2282.get(0);
        mod_2281.put(0, t);
    endrule
    rule rule_2947;
        ChannelMessage t;
        t <- mod_2271.get(0);
        mod_2273.put(0, t);
    endrule
    rule rule_2948;
        ChannelMessage t;
        t <- mod_2271.get(1);
        mod_2272.put(1, t);
    endrule
    rule rule_2949;
        ChannelMessage t;
        t <- mod_2281.get(0);
        mod_2280.put(0, t);
    endrule
    rule rule_2950;
        ChannelMessage t;
        t <- mod_2284.get(0);
        mod_2283.put(1, t);
    endrule
    rule rule_2951;
        ChannelMessage t;
        t <- mod_2267.get(0);
        mod_2279.put(0, t);
    endrule
    rule rule_2952;
        ChannelMessage t;
        t <- mod_2273.get(0);
        mod_2273.put(1, t);
    endrule
    rule rule_2953;
        ChannelMessage t;
        t <- mod_2267.get(1);
        mod_2268.put(0, t);
    endrule
    rule rule_2954;
        ChannelMessage t;
        t <- mod_2261.get(1);
        mod_2262.put(0, t);
    endrule
    rule rule_2955;
        ChannelMessage t;
        t <- mod_2261.get(0);
        mod_2294.put(0, t);
    endrule
    rule rule_2956;
        ChannelMessage t;
        t <- mod_2263.get(1);
        mod_2264.put(0, t);
    endrule
    rule rule_2957;
        ChannelMessage t;
        t <- mod_2260.get(3);
        mod_2261.put(0, t);
    endrule
    rule rule_2958;
        ChannelMessage t;
        t <- mod_2275.get(0);
        mod_2276.put(0, t);
    endrule
    rule rule_2959;
        ChannelMessage t;
        t <- mod_2274.get(1);
        mod_2270.put(1, t);
    endrule
    rule rule_2960;
        ChannelMessage t;
        t <- mod_2279.get(0);
        mod_2267.put(1, t);
    endrule
    rule rule_2961;
        ChannelMessage t;
        t <- mod_2285.get(0);
        mod_2283.put(0, t);
    endrule
    rule rule_2962;
        ChannelMessage t;
        t <- mod_2289.get(0);
        mod_2290.put(0, t);
    endrule
    rule rule_2963;
        ChannelMessage t;
        t <- mod_2275.get(1);
        mod_2268.put(1, t);
    endrule
    rule rule_2964;
        ChannelMessage t;
        t <- mod_2288.get(0);
        mod_2287.put(1, t);
    endrule
    rule rule_2965;
        ChannelMessage t;
        t <- mod_2265.get(0);
        mod_2266.put(0, t);
    endrule
    rule rule_2966;
        ChannelMessage t;
        t <- mod_2277.get(0);
        mod_2275.put(0, t);
    endrule
    rule rule_2967;
        ChannelMessage t;
        t <- mod_2262.get(1);
        mod_2263.put(0, t);
    endrule
    rule rule_2968;
        ChannelMessage t;
        t <- mod_2258.get(0);
        mod_2259.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2256.put(0, t);
        end
        if (i == 1) begin
            mod_2272.put(0, t);
        end
        if (i == 2) begin
            mod_2278.put(0, t);
        end
        if (i == 3) begin
            mod_2286.put(0, t);
        end
        if (i == 4) begin
            mod_2292.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_2260.get(0);
        end
        if (i == 1) begin
            t <- mod_2260.get(1);
        end
        if (i == 3) begin
            t <- mod_2260.get(2);
        end
        if (i == 2) begin
            t <- mod_2272.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6090 (Operation_IFC);
    Operation_IFC mod_2297_inner <- mkReshape(2, 64);
    Operation_IFC mod_2297 <- mkDebugOperation(mod_2297_inner, "mod_2297");
    Operation_IFC mod_2298_inner <- mkFlatten(1);
    Operation_IFC mod_2298 <- mkDebugOperation(mod_2298_inner, "mod_2298");
    Operation_IFC mod_2299_inner <- mkFlatten(2);
    Operation_IFC mod_2299 <- mkDebugOperation(mod_2299_inner, "mod_2299");
    Operation_IFC mod_2300_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2300 <- mkDebugOperation(mod_2300_inner, "mod_2300");
    Broadcast_IFC#(4) mod_2301_inner <- mkBroadcast(4);
    Operation_IFC mod_2301 <- mkDebugOperation(mod_2301_inner.op, "mod_2301");
    PMU_IFC mod_2302_bufferize <- mkPMU(2);
    Operation_IFC mod_2302_inner = mod_2302_bufferize.operation;
    Operation_IFC mod_2302 <- mkDebugOperation(mod_2302_inner, "mod_2302");
    Broadcast_IFC#(2) mod_2303_inner <- mkBroadcast(2);
    Operation_IFC mod_2303 <- mkDebugOperation(mod_2303_inner.op, "mod_2303");
    PMU_IFC mod_2304_bufferize <- mkPMU(1);
    Operation_IFC mod_2304_inner = mod_2304_bufferize.operation;
    Operation_IFC mod_2304 <- mkDebugOperation(mod_2304_inner, "mod_2304");
    Operation_IFC mod_2305_inner <- mkBinaryMap(1100, matmul_t_tile);
    Operation_IFC mod_2305 <- mkDebugOperation(mod_2305_inner, "mod_2305");
    Operation_IFC mod_2306_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2306 <- mkDebugOperation(mod_2306_inner, "mod_2306");
    Operation_IFC mod_2307_inner <- mkBinaryMap(1868, mul_tile);
    Operation_IFC mod_2307 <- mkDebugOperation(mod_2307_inner, "mod_2307");
    PMU_IFC mod_2308_bufferize <- mkPMU(1);
    Operation_IFC mod_2308_inner = mod_2308_bufferize.operation;
    Operation_IFC mod_2308 <- mkDebugOperation(mod_2308_inner, "mod_2308");
    Operation_IFC mod_2309_inner <- mkBinaryMap(2451, matmul_t_tile);
    Operation_IFC mod_2309 <- mkDebugOperation(mod_2309_inner, "mod_2309");
    Operation_IFC mod_2310_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2310 <- mkDebugOperation(mod_2310_inner, "mod_2310");
    Operation_IFC mod_2311_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2311 <- mkDebugOperation(mod_2311_inner, "mod_2311");
    Operation_IFC mod_2312_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2312 <- mkDebugOperation(mod_2312_inner, "mod_2312");
    Operation_IFC mod_2313_inner <- mkBinaryMap(2767, mul_tile);
    Operation_IFC mod_2313 <- mkDebugOperation(mod_2313_inner, "mod_2313");
    PMU_IFC mod_2314_bufferize <- mkPMU(1);
    Operation_IFC mod_2314_inner = mod_2314_bufferize.operation;
    Operation_IFC mod_2314 <- mkDebugOperation(mod_2314_inner, "mod_2314");
    PMU_IFC mod_2315_bufferize <- mkPMU(2);
    Operation_IFC mod_2315_inner = mod_2315_bufferize.operation;
    Operation_IFC mod_2315 <- mkDebugOperation(mod_2315_inner, "mod_2315");
    PMU_IFC mod_2316_bufferize <- mkPMU(2);
    Operation_IFC mod_2316_inner = mod_2316_bufferize.operation;
    Operation_IFC mod_2316 <- mkDebugOperation(mod_2316_inner, "mod_2316");
    Operation_IFC mod_2317_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2317 <- mkDebugOperation(mod_2317_inner, "mod_2317");
    Operation_IFC mod_2318_inner <- mkFlatten(1);
    Operation_IFC mod_2318 <- mkDebugOperation(mod_2318_inner, "mod_2318");
    Operation_IFC mod_2319_inner <- mkFlatten(0);
    Operation_IFC mod_2319 <- mkDebugOperation(mod_2319_inner, "mod_2319");
    Operation_IFC mod_2320_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2320 <- mkDebugOperation(mod_2320_inner, "mod_2320");
    Operation_IFC mod_2321_inner <- mkUnaryMap(1740, silu_tile);
    Operation_IFC mod_2321 <- mkDebugOperation(mod_2321_inner, "mod_2321");
    Operation_IFC mod_2322_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2322 <- mkDebugOperation(mod_2322_inner, "mod_2322");
    Operation_IFC mod_2323_inner <- mkBinaryMap(1612, matmul_t_tile);
    Operation_IFC mod_2323 <- mkDebugOperation(mod_2323_inner, "mod_2323");
    PMU_IFC mod_2324_bufferize <- mkPMU(2);
    Operation_IFC mod_2324_inner = mod_2324_bufferize.operation;
    Operation_IFC mod_2324 <- mkDebugOperation(mod_2324_inner, "mod_2324");
    Operation_IFC mod_2325_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2325 <- mkDebugOperation(mod_2325_inner, "mod_2325");
    Operation_IFC mod_2326_inner <- mkFlatten(1);
    Operation_IFC mod_2326 <- mkDebugOperation(mod_2326_inner, "mod_2326");
    Operation_IFC mod_2327_inner <- mkFlatten(0);
    Operation_IFC mod_2327 <- mkDebugOperation(mod_2327_inner, "mod_2327");
    PMU_IFC mod_2328_bufferize <- mkPMU(1);
    Operation_IFC mod_2328_inner = mod_2328_bufferize.operation;
    Operation_IFC mod_2328 <- mkDebugOperation(mod_2328_inner, "mod_2328");
    Operation_IFC mod_2329_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2329 <- mkDebugOperation(mod_2329_inner, "mod_2329");
    PMU_IFC mod_2330_bufferize <- mkPMU(2);
    Operation_IFC mod_2330_inner = mod_2330_bufferize.operation;
    Operation_IFC mod_2330 <- mkDebugOperation(mod_2330_inner, "mod_2330");
    Operation_IFC mod_2331_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2331 <- mkDebugOperation(mod_2331_inner, "mod_2331");
    Operation_IFC mod_2332_inner <- mkFlatten(1);
    Operation_IFC mod_2332 <- mkDebugOperation(mod_2332_inner, "mod_2332");
    Operation_IFC mod_2333_inner <- mkFlatten(0);
    Operation_IFC mod_2333 <- mkDebugOperation(mod_2333_inner, "mod_2333");
    Operation_IFC mod_2334_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2334 <- mkDebugOperation(mod_2334_inner, "mod_2334");
    Operation_IFC mod_2335_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2335 <- mkDebugOperation(mod_2335_inner, "mod_2335");
    PMU_IFC mod_2336_bufferize <- mkPMU(2);
    Operation_IFC mod_2336_inner = mod_2336_bufferize.operation;
    Operation_IFC mod_2336 <- mkDebugOperation(mod_2336_inner, "mod_2336");
    rule rule_2969;
        ChannelMessage t;
        t <- mod_2325.get(0);
        mod_2324.put(1, t);
    endrule
    rule rule_2970;
        ChannelMessage t;
        t <- mod_2329.get(0);
        mod_2328.put(1, t);
    endrule
    rule rule_2971;
        ChannelMessage t;
        t <- mod_2311.get(1);
        mod_2312.put(0, t);
    endrule
    rule rule_2972;
        ChannelMessage t;
        t <- mod_2303.get(1);
        mod_2304.put(0, t);
    endrule
    rule rule_2973;
        ChannelMessage t;
        t <- mod_2312.get(0);
        mod_2314.put(0, t);
    endrule
    rule rule_2974;
        ChannelMessage t;
        t <- mod_2321.get(0);
        mod_2307.put(1, t);
    endrule
    rule rule_2975;
        ChannelMessage t;
        t <- mod_2335.get(0);
        mod_2302.put(1, t);
    endrule
    rule rule_2976;
        ChannelMessage t;
        t <- mod_2336.get(0);
        mod_2336.put(1, t);
    endrule
    rule rule_2977;
        ChannelMessage t;
        t <- mod_2324.get(1);
        mod_2323.put(1, t);
    endrule
    rule rule_2978;
        ChannelMessage t;
        t <- mod_2328.get(0);
        mod_2329.put(0, t);
    endrule
    rule rule_2979;
        ChannelMessage t;
        t <- mod_2315.get(1);
        mod_2311.put(1, t);
    endrule
    rule rule_2980;
        ChannelMessage t;
        t <- mod_2331.get(0);
        mod_2330.put(1, t);
    endrule
    rule rule_2981;
        ChannelMessage t;
        t <- mod_2318.get(0);
        mod_2316.put(0, t);
    endrule
    rule rule_2982;
        ChannelMessage t;
        t <- mod_2305.get(0);
        mod_2306.put(0, t);
    endrule
    rule rule_2983;
        ChannelMessage t;
        t <- mod_2311.get(0);
        mod_2315.put(0, t);
    endrule
    rule rule_2984;
        ChannelMessage t;
        t <- mod_2323.get(0);
        mod_2322.put(0, t);
    endrule
    rule rule_2985;
        ChannelMessage t;
        t <- mod_2322.get(0);
        mod_2321.put(0, t);
    endrule
    rule rule_2986;
        ChannelMessage t;
        t <- mod_2336.get(1);
        mod_2300.put(1, t);
    endrule
    rule rule_2987;
        ChannelMessage t;
        t <- mod_2332.get(0);
        mod_2330.put(0, t);
    endrule
    rule rule_2988;
        ChannelMessage t;
        t <- mod_2326.get(0);
        mod_2324.put(0, t);
    endrule
    rule rule_2989;
        ChannelMessage t;
        t <- mod_2316.get(0);
        mod_2317.put(0, t);
    endrule
    rule rule_2990;
        ChannelMessage t;
        t <- mod_2314.get(1);
        mod_2312.put(1, t);
    endrule
    rule rule_2991;
        ChannelMessage t;
        t <- mod_2300.get(0);
        mod_2336.put(0, t);
    endrule
    rule rule_2992;
        ChannelMessage t;
        t <- mod_2298.get(0);
        mod_2299.put(0, t);
    endrule
    rule rule_2993;
        ChannelMessage t;
        t <- mod_2319.get(0);
        mod_2318.put(0, t);
    endrule
    rule rule_2994;
        ChannelMessage t;
        t <- mod_2324.get(0);
        mod_2325.put(0, t);
    endrule
    rule rule_2995;
        ChannelMessage t;
        t <- mod_2327.get(0);
        mod_2326.put(0, t);
    endrule
    rule rule_2996;
        ChannelMessage t;
        t <- mod_2300.get(1);
        mod_2301.put(0, t);
    endrule
    rule rule_2997;
        ChannelMessage t;
        t <- mod_2328.get(1);
        mod_2323.put(0, t);
    endrule
    rule rule_2998;
        ChannelMessage t;
        t <- mod_2304.get(1);
        mod_2305.put(0, t);
    endrule
    rule rule_2999;
        ChannelMessage t;
        t <- mod_2309.get(0);
        mod_2310.put(0, t);
    endrule
    rule rule_3000;
        ChannelMessage t;
        t <- mod_2308.get(0);
        mod_2320.put(0, t);
    endrule
    rule rule_3001;
        ChannelMessage t;
        t <- mod_2308.get(1);
        mod_2309.put(0, t);
    endrule
    rule rule_3002;
        ChannelMessage t;
        t <- mod_2320.get(0);
        mod_2308.put(1, t);
    endrule
    rule rule_3003;
        ChannelMessage t;
        t <- mod_2297.get(0);
        mod_2298.put(0, t);
    endrule
    rule rule_3004;
        ChannelMessage t;
        t <- mod_2312.get(1);
        mod_2313.put(1, t);
    endrule
    rule rule_3005;
        ChannelMessage t;
        t <- mod_2330.get(0);
        mod_2331.put(0, t);
    endrule
    rule rule_3006;
        ChannelMessage t;
        t <- mod_2315.get(0);
        mod_2315.put(1, t);
    endrule
    rule rule_3007;
        ChannelMessage t;
        t <- mod_2307.get(0);
        mod_2308.put(0, t);
    endrule
    rule rule_3008;
        ChannelMessage t;
        t <- mod_2301.get(3);
        mod_2302.put(0, t);
    endrule
    rule rule_3009;
        ChannelMessage t;
        t <- mod_2333.get(0);
        mod_2332.put(0, t);
    endrule
    rule rule_3010;
        ChannelMessage t;
        t <- mod_2316.get(1);
        mod_2309.put(1, t);
    endrule
    rule rule_3011;
        ChannelMessage t;
        t <- mod_2302.get(0);
        mod_2335.put(0, t);
    endrule
    rule rule_3012;
        ChannelMessage t;
        t <- mod_2304.get(0);
        mod_2334.put(0, t);
    endrule
    rule rule_3013;
        ChannelMessage t;
        t <- mod_2306.get(0);
        mod_2307.put(0, t);
    endrule
    rule rule_3014;
        ChannelMessage t;
        t <- mod_2302.get(1);
        mod_2303.put(0, t);
    endrule
    rule rule_3015;
        ChannelMessage t;
        t <- mod_2310.get(0);
        mod_2311.put(0, t);
    endrule
    rule rule_3016;
        ChannelMessage t;
        t <- mod_2317.get(0);
        mod_2316.put(1, t);
    endrule
    rule rule_3017;
        ChannelMessage t;
        t <- mod_2334.get(0);
        mod_2304.put(1, t);
    endrule
    rule rule_3018;
        ChannelMessage t;
        t <- mod_2299.get(0);
        mod_2300.put(0, t);
    endrule
    rule rule_3019;
        ChannelMessage t;
        t <- mod_2330.get(1);
        mod_2305.put(1, t);
    endrule
    rule rule_3020;
        ChannelMessage t;
        t <- mod_2314.get(0);
        mod_2314.put(1, t);
    endrule
    rule rule_3021;
        ChannelMessage t;
        t <- mod_2303.get(0);
        mod_2328.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2297.put(0, t);
        end
        if (i == 1) begin
            mod_2313.put(0, t);
        end
        if (i == 2) begin
            mod_2319.put(0, t);
        end
        if (i == 3) begin
            mod_2327.put(0, t);
        end
        if (i == 4) begin
            mod_2333.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 2) begin
            t <- mod_2301.get(0);
        end
        if (i == 3) begin
            t <- mod_2301.get(1);
        end
        if (i == 0) begin
            t <- mod_2301.get(2);
        end
        if (i == 1) begin
            t <- mod_2313.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6091 (Operation_IFC);
    Operation_IFC mod_2338_inner <- mkReshape(2, 64);
    Operation_IFC mod_2338 <- mkDebugOperation(mod_2338_inner, "mod_2338");
    Operation_IFC mod_2339_inner <- mkFlatten(1);
    Operation_IFC mod_2339 <- mkDebugOperation(mod_2339_inner, "mod_2339");
    Operation_IFC mod_2340_inner <- mkFlatten(2);
    Operation_IFC mod_2340 <- mkDebugOperation(mod_2340_inner, "mod_2340");
    Operation_IFC mod_2341_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2341 <- mkDebugOperation(mod_2341_inner, "mod_2341");
    Broadcast_IFC#(4) mod_2342_inner <- mkBroadcast(4);
    Operation_IFC mod_2342 <- mkDebugOperation(mod_2342_inner.op, "mod_2342");
    PMU_IFC mod_2343_bufferize <- mkPMU(2);
    Operation_IFC mod_2343_inner = mod_2343_bufferize.operation;
    Operation_IFC mod_2343 <- mkDebugOperation(mod_2343_inner, "mod_2343");
    Broadcast_IFC#(2) mod_2344_inner <- mkBroadcast(2);
    Operation_IFC mod_2344 <- mkDebugOperation(mod_2344_inner.op, "mod_2344");
    PMU_IFC mod_2345_bufferize <- mkPMU(1);
    Operation_IFC mod_2345_inner = mod_2345_bufferize.operation;
    Operation_IFC mod_2345 <- mkDebugOperation(mod_2345_inner, "mod_2345");
    Operation_IFC mod_2346_inner <- mkBinaryMap(1099, matmul_t_tile);
    Operation_IFC mod_2346 <- mkDebugOperation(mod_2346_inner, "mod_2346");
    Operation_IFC mod_2347_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2347 <- mkDebugOperation(mod_2347_inner, "mod_2347");
    Operation_IFC mod_2348_inner <- mkBinaryMap(1867, mul_tile);
    Operation_IFC mod_2348 <- mkDebugOperation(mod_2348_inner, "mod_2348");
    PMU_IFC mod_2349_bufferize <- mkPMU(1);
    Operation_IFC mod_2349_inner = mod_2349_bufferize.operation;
    Operation_IFC mod_2349 <- mkDebugOperation(mod_2349_inner, "mod_2349");
    Operation_IFC mod_2350_inner <- mkBinaryMap(2449, matmul_t_tile);
    Operation_IFC mod_2350 <- mkDebugOperation(mod_2350_inner, "mod_2350");
    Operation_IFC mod_2351_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2351 <- mkDebugOperation(mod_2351_inner, "mod_2351");
    Operation_IFC mod_2352_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2352 <- mkDebugOperation(mod_2352_inner, "mod_2352");
    Operation_IFC mod_2353_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2353 <- mkDebugOperation(mod_2353_inner, "mod_2353");
    Operation_IFC mod_2354_inner <- mkBinaryMap(2766, mul_tile);
    Operation_IFC mod_2354 <- mkDebugOperation(mod_2354_inner, "mod_2354");
    PMU_IFC mod_2355_bufferize <- mkPMU(1);
    Operation_IFC mod_2355_inner = mod_2355_bufferize.operation;
    Operation_IFC mod_2355 <- mkDebugOperation(mod_2355_inner, "mod_2355");
    PMU_IFC mod_2356_bufferize <- mkPMU(2);
    Operation_IFC mod_2356_inner = mod_2356_bufferize.operation;
    Operation_IFC mod_2356 <- mkDebugOperation(mod_2356_inner, "mod_2356");
    PMU_IFC mod_2357_bufferize <- mkPMU(2);
    Operation_IFC mod_2357_inner = mod_2357_bufferize.operation;
    Operation_IFC mod_2357 <- mkDebugOperation(mod_2357_inner, "mod_2357");
    Operation_IFC mod_2358_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2358 <- mkDebugOperation(mod_2358_inner, "mod_2358");
    Operation_IFC mod_2359_inner <- mkFlatten(1);
    Operation_IFC mod_2359 <- mkDebugOperation(mod_2359_inner, "mod_2359");
    Operation_IFC mod_2360_inner <- mkFlatten(0);
    Operation_IFC mod_2360 <- mkDebugOperation(mod_2360_inner, "mod_2360");
    Operation_IFC mod_2361_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2361 <- mkDebugOperation(mod_2361_inner, "mod_2361");
    Operation_IFC mod_2362_inner <- mkUnaryMap(1739, silu_tile);
    Operation_IFC mod_2362 <- mkDebugOperation(mod_2362_inner, "mod_2362");
    Operation_IFC mod_2363_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2363 <- mkDebugOperation(mod_2363_inner, "mod_2363");
    Operation_IFC mod_2364_inner <- mkBinaryMap(1611, matmul_t_tile);
    Operation_IFC mod_2364 <- mkDebugOperation(mod_2364_inner, "mod_2364");
    PMU_IFC mod_2365_bufferize <- mkPMU(2);
    Operation_IFC mod_2365_inner = mod_2365_bufferize.operation;
    Operation_IFC mod_2365 <- mkDebugOperation(mod_2365_inner, "mod_2365");
    Operation_IFC mod_2366_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2366 <- mkDebugOperation(mod_2366_inner, "mod_2366");
    Operation_IFC mod_2367_inner <- mkFlatten(1);
    Operation_IFC mod_2367 <- mkDebugOperation(mod_2367_inner, "mod_2367");
    Operation_IFC mod_2368_inner <- mkFlatten(0);
    Operation_IFC mod_2368 <- mkDebugOperation(mod_2368_inner, "mod_2368");
    PMU_IFC mod_2369_bufferize <- mkPMU(1);
    Operation_IFC mod_2369_inner = mod_2369_bufferize.operation;
    Operation_IFC mod_2369 <- mkDebugOperation(mod_2369_inner, "mod_2369");
    Operation_IFC mod_2370_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2370 <- mkDebugOperation(mod_2370_inner, "mod_2370");
    PMU_IFC mod_2371_bufferize <- mkPMU(2);
    Operation_IFC mod_2371_inner = mod_2371_bufferize.operation;
    Operation_IFC mod_2371 <- mkDebugOperation(mod_2371_inner, "mod_2371");
    Operation_IFC mod_2372_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2372 <- mkDebugOperation(mod_2372_inner, "mod_2372");
    Operation_IFC mod_2373_inner <- mkFlatten(1);
    Operation_IFC mod_2373 <- mkDebugOperation(mod_2373_inner, "mod_2373");
    Operation_IFC mod_2374_inner <- mkFlatten(0);
    Operation_IFC mod_2374 <- mkDebugOperation(mod_2374_inner, "mod_2374");
    Operation_IFC mod_2375_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2375 <- mkDebugOperation(mod_2375_inner, "mod_2375");
    Operation_IFC mod_2376_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2376 <- mkDebugOperation(mod_2376_inner, "mod_2376");
    PMU_IFC mod_2377_bufferize <- mkPMU(2);
    Operation_IFC mod_2377_inner = mod_2377_bufferize.operation;
    Operation_IFC mod_2377 <- mkDebugOperation(mod_2377_inner, "mod_2377");
    rule rule_3022;
        ChannelMessage t;
        t <- mod_2343.get(1);
        mod_2344.put(0, t);
    endrule
    rule rule_3023;
        ChannelMessage t;
        t <- mod_2344.get(1);
        mod_2345.put(0, t);
    endrule
    rule rule_3024;
        ChannelMessage t;
        t <- mod_2375.get(0);
        mod_2345.put(1, t);
    endrule
    rule rule_3025;
        ChannelMessage t;
        t <- mod_2347.get(0);
        mod_2348.put(0, t);
    endrule
    rule rule_3026;
        ChannelMessage t;
        t <- mod_2350.get(0);
        mod_2351.put(0, t);
    endrule
    rule rule_3027;
        ChannelMessage t;
        t <- mod_2351.get(0);
        mod_2352.put(0, t);
    endrule
    rule rule_3028;
        ChannelMessage t;
        t <- mod_2349.get(1);
        mod_2350.put(0, t);
    endrule
    rule rule_3029;
        ChannelMessage t;
        t <- mod_2353.get(0);
        mod_2355.put(0, t);
    endrule
    rule rule_3030;
        ChannelMessage t;
        t <- mod_2348.get(0);
        mod_2349.put(0, t);
    endrule
    rule rule_3031;
        ChannelMessage t;
        t <- mod_2369.get(1);
        mod_2364.put(0, t);
    endrule
    rule rule_3032;
        ChannelMessage t;
        t <- mod_2340.get(0);
        mod_2341.put(0, t);
    endrule
    rule rule_3033;
        ChannelMessage t;
        t <- mod_2338.get(0);
        mod_2339.put(0, t);
    endrule
    rule rule_3034;
        ChannelMessage t;
        t <- mod_2346.get(0);
        mod_2347.put(0, t);
    endrule
    rule rule_3035;
        ChannelMessage t;
        t <- mod_2377.get(1);
        mod_2341.put(1, t);
    endrule
    rule rule_3036;
        ChannelMessage t;
        t <- mod_2352.get(1);
        mod_2353.put(0, t);
    endrule
    rule rule_3037;
        ChannelMessage t;
        t <- mod_2377.get(0);
        mod_2377.put(1, t);
    endrule
    rule rule_3038;
        ChannelMessage t;
        t <- mod_2374.get(0);
        mod_2373.put(0, t);
    endrule
    rule rule_3039;
        ChannelMessage t;
        t <- mod_2356.get(1);
        mod_2352.put(1, t);
    endrule
    rule rule_3040;
        ChannelMessage t;
        t <- mod_2366.get(0);
        mod_2365.put(1, t);
    endrule
    rule rule_3041;
        ChannelMessage t;
        t <- mod_2355.get(1);
        mod_2353.put(1, t);
    endrule
    rule rule_3042;
        ChannelMessage t;
        t <- mod_2361.get(0);
        mod_2349.put(1, t);
    endrule
    rule rule_3043;
        ChannelMessage t;
        t <- mod_2367.get(0);
        mod_2365.put(0, t);
    endrule
    rule rule_3044;
        ChannelMessage t;
        t <- mod_2341.get(0);
        mod_2377.put(0, t);
    endrule
    rule rule_3045;
        ChannelMessage t;
        t <- mod_2339.get(0);
        mod_2340.put(0, t);
    endrule
    rule rule_3046;
        ChannelMessage t;
        t <- mod_2353.get(1);
        mod_2354.put(1, t);
    endrule
    rule rule_3047;
        ChannelMessage t;
        t <- mod_2363.get(0);
        mod_2362.put(0, t);
    endrule
    rule rule_3048;
        ChannelMessage t;
        t <- mod_2343.get(0);
        mod_2376.put(0, t);
    endrule
    rule rule_3049;
        ChannelMessage t;
        t <- mod_2349.get(0);
        mod_2361.put(0, t);
    endrule
    rule rule_3050;
        ChannelMessage t;
        t <- mod_2345.get(1);
        mod_2346.put(0, t);
    endrule
    rule rule_3051;
        ChannelMessage t;
        t <- mod_2360.get(0);
        mod_2359.put(0, t);
    endrule
    rule rule_3052;
        ChannelMessage t;
        t <- mod_2362.get(0);
        mod_2348.put(1, t);
    endrule
    rule rule_3053;
        ChannelMessage t;
        t <- mod_2371.get(1);
        mod_2346.put(1, t);
    endrule
    rule rule_3054;
        ChannelMessage t;
        t <- mod_2355.get(0);
        mod_2355.put(1, t);
    endrule
    rule rule_3055;
        ChannelMessage t;
        t <- mod_2341.get(1);
        mod_2342.put(0, t);
    endrule
    rule rule_3056;
        ChannelMessage t;
        t <- mod_2370.get(0);
        mod_2369.put(1, t);
    endrule
    rule rule_3057;
        ChannelMessage t;
        t <- mod_2364.get(0);
        mod_2363.put(0, t);
    endrule
    rule rule_3058;
        ChannelMessage t;
        t <- mod_2371.get(0);
        mod_2372.put(0, t);
    endrule
    rule rule_3059;
        ChannelMessage t;
        t <- mod_2373.get(0);
        mod_2371.put(0, t);
    endrule
    rule rule_3060;
        ChannelMessage t;
        t <- mod_2342.get(3);
        mod_2343.put(0, t);
    endrule
    rule rule_3061;
        ChannelMessage t;
        t <- mod_2358.get(0);
        mod_2357.put(1, t);
    endrule
    rule rule_3062;
        ChannelMessage t;
        t <- mod_2369.get(0);
        mod_2370.put(0, t);
    endrule
    rule rule_3063;
        ChannelMessage t;
        t <- mod_2357.get(0);
        mod_2358.put(0, t);
    endrule
    rule rule_3064;
        ChannelMessage t;
        t <- mod_2357.get(1);
        mod_2350.put(1, t);
    endrule
    rule rule_3065;
        ChannelMessage t;
        t <- mod_2345.get(0);
        mod_2375.put(0, t);
    endrule
    rule rule_3066;
        ChannelMessage t;
        t <- mod_2376.get(0);
        mod_2343.put(1, t);
    endrule
    rule rule_3067;
        ChannelMessage t;
        t <- mod_2352.get(0);
        mod_2356.put(0, t);
    endrule
    rule rule_3068;
        ChannelMessage t;
        t <- mod_2365.get(0);
        mod_2366.put(0, t);
    endrule
    rule rule_3069;
        ChannelMessage t;
        t <- mod_2368.get(0);
        mod_2367.put(0, t);
    endrule
    rule rule_3070;
        ChannelMessage t;
        t <- mod_2344.get(0);
        mod_2369.put(0, t);
    endrule
    rule rule_3071;
        ChannelMessage t;
        t <- mod_2365.get(1);
        mod_2364.put(1, t);
    endrule
    rule rule_3072;
        ChannelMessage t;
        t <- mod_2372.get(0);
        mod_2371.put(1, t);
    endrule
    rule rule_3073;
        ChannelMessage t;
        t <- mod_2356.get(0);
        mod_2356.put(1, t);
    endrule
    rule rule_3074;
        ChannelMessage t;
        t <- mod_2359.get(0);
        mod_2357.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2338.put(0, t);
        end
        if (i == 1) begin
            mod_2354.put(0, t);
        end
        if (i == 2) begin
            mod_2360.put(0, t);
        end
        if (i == 3) begin
            mod_2368.put(0, t);
        end
        if (i == 4) begin
            mod_2374.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_2342.get(0);
        end
        if (i == 2) begin
            t <- mod_2342.get(1);
        end
        if (i == 0) begin
            t <- mod_2342.get(2);
        end
        if (i == 1) begin
            t <- mod_2354.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6092 (Operation_IFC);
    Operation_IFC mod_2379_inner <- mkReshape(2, 64);
    Operation_IFC mod_2379 <- mkDebugOperation(mod_2379_inner, "mod_2379");
    Operation_IFC mod_2380_inner <- mkFlatten(1);
    Operation_IFC mod_2380 <- mkDebugOperation(mod_2380_inner, "mod_2380");
    Operation_IFC mod_2381_inner <- mkFlatten(2);
    Operation_IFC mod_2381 <- mkDebugOperation(mod_2381_inner, "mod_2381");
    Operation_IFC mod_2382_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2382 <- mkDebugOperation(mod_2382_inner, "mod_2382");
    Broadcast_IFC#(4) mod_2383_inner <- mkBroadcast(4);
    Operation_IFC mod_2383 <- mkDebugOperation(mod_2383_inner.op, "mod_2383");
    PMU_IFC mod_2384_bufferize <- mkPMU(2);
    Operation_IFC mod_2384_inner = mod_2384_bufferize.operation;
    Operation_IFC mod_2384 <- mkDebugOperation(mod_2384_inner, "mod_2384");
    Broadcast_IFC#(2) mod_2385_inner <- mkBroadcast(2);
    Operation_IFC mod_2385 <- mkDebugOperation(mod_2385_inner.op, "mod_2385");
    PMU_IFC mod_2386_bufferize <- mkPMU(1);
    Operation_IFC mod_2386_inner = mod_2386_bufferize.operation;
    Operation_IFC mod_2386 <- mkDebugOperation(mod_2386_inner, "mod_2386");
    Operation_IFC mod_2387_inner <- mkBinaryMap(1098, matmul_t_tile);
    Operation_IFC mod_2387 <- mkDebugOperation(mod_2387_inner, "mod_2387");
    Operation_IFC mod_2388_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2388 <- mkDebugOperation(mod_2388_inner, "mod_2388");
    Operation_IFC mod_2389_inner <- mkBinaryMap(1866, mul_tile);
    Operation_IFC mod_2389 <- mkDebugOperation(mod_2389_inner, "mod_2389");
    PMU_IFC mod_2390_bufferize <- mkPMU(1);
    Operation_IFC mod_2390_inner = mod_2390_bufferize.operation;
    Operation_IFC mod_2390 <- mkDebugOperation(mod_2390_inner, "mod_2390");
    Operation_IFC mod_2391_inner <- mkBinaryMap(2447, matmul_t_tile);
    Operation_IFC mod_2391 <- mkDebugOperation(mod_2391_inner, "mod_2391");
    Operation_IFC mod_2392_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2392 <- mkDebugOperation(mod_2392_inner, "mod_2392");
    Operation_IFC mod_2393_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2393 <- mkDebugOperation(mod_2393_inner, "mod_2393");
    Operation_IFC mod_2394_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2394 <- mkDebugOperation(mod_2394_inner, "mod_2394");
    Operation_IFC mod_2395_inner <- mkBinaryMap(2765, mul_tile);
    Operation_IFC mod_2395 <- mkDebugOperation(mod_2395_inner, "mod_2395");
    PMU_IFC mod_2396_bufferize <- mkPMU(1);
    Operation_IFC mod_2396_inner = mod_2396_bufferize.operation;
    Operation_IFC mod_2396 <- mkDebugOperation(mod_2396_inner, "mod_2396");
    PMU_IFC mod_2397_bufferize <- mkPMU(2);
    Operation_IFC mod_2397_inner = mod_2397_bufferize.operation;
    Operation_IFC mod_2397 <- mkDebugOperation(mod_2397_inner, "mod_2397");
    PMU_IFC mod_2398_bufferize <- mkPMU(2);
    Operation_IFC mod_2398_inner = mod_2398_bufferize.operation;
    Operation_IFC mod_2398 <- mkDebugOperation(mod_2398_inner, "mod_2398");
    Operation_IFC mod_2399_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2399 <- mkDebugOperation(mod_2399_inner, "mod_2399");
    Operation_IFC mod_2400_inner <- mkFlatten(1);
    Operation_IFC mod_2400 <- mkDebugOperation(mod_2400_inner, "mod_2400");
    Operation_IFC mod_2401_inner <- mkFlatten(0);
    Operation_IFC mod_2401 <- mkDebugOperation(mod_2401_inner, "mod_2401");
    Operation_IFC mod_2402_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2402 <- mkDebugOperation(mod_2402_inner, "mod_2402");
    Operation_IFC mod_2403_inner <- mkUnaryMap(1738, silu_tile);
    Operation_IFC mod_2403 <- mkDebugOperation(mod_2403_inner, "mod_2403");
    Operation_IFC mod_2404_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2404 <- mkDebugOperation(mod_2404_inner, "mod_2404");
    Operation_IFC mod_2405_inner <- mkBinaryMap(1610, matmul_t_tile);
    Operation_IFC mod_2405 <- mkDebugOperation(mod_2405_inner, "mod_2405");
    PMU_IFC mod_2406_bufferize <- mkPMU(2);
    Operation_IFC mod_2406_inner = mod_2406_bufferize.operation;
    Operation_IFC mod_2406 <- mkDebugOperation(mod_2406_inner, "mod_2406");
    Operation_IFC mod_2407_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2407 <- mkDebugOperation(mod_2407_inner, "mod_2407");
    Operation_IFC mod_2408_inner <- mkFlatten(1);
    Operation_IFC mod_2408 <- mkDebugOperation(mod_2408_inner, "mod_2408");
    Operation_IFC mod_2409_inner <- mkFlatten(0);
    Operation_IFC mod_2409 <- mkDebugOperation(mod_2409_inner, "mod_2409");
    PMU_IFC mod_2410_bufferize <- mkPMU(1);
    Operation_IFC mod_2410_inner = mod_2410_bufferize.operation;
    Operation_IFC mod_2410 <- mkDebugOperation(mod_2410_inner, "mod_2410");
    Operation_IFC mod_2411_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2411 <- mkDebugOperation(mod_2411_inner, "mod_2411");
    PMU_IFC mod_2412_bufferize <- mkPMU(2);
    Operation_IFC mod_2412_inner = mod_2412_bufferize.operation;
    Operation_IFC mod_2412 <- mkDebugOperation(mod_2412_inner, "mod_2412");
    Operation_IFC mod_2413_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2413 <- mkDebugOperation(mod_2413_inner, "mod_2413");
    Operation_IFC mod_2414_inner <- mkFlatten(1);
    Operation_IFC mod_2414 <- mkDebugOperation(mod_2414_inner, "mod_2414");
    Operation_IFC mod_2415_inner <- mkFlatten(0);
    Operation_IFC mod_2415 <- mkDebugOperation(mod_2415_inner, "mod_2415");
    Operation_IFC mod_2416_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2416 <- mkDebugOperation(mod_2416_inner, "mod_2416");
    Operation_IFC mod_2417_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2417 <- mkDebugOperation(mod_2417_inner, "mod_2417");
    PMU_IFC mod_2418_bufferize <- mkPMU(2);
    Operation_IFC mod_2418_inner = mod_2418_bufferize.operation;
    Operation_IFC mod_2418 <- mkDebugOperation(mod_2418_inner, "mod_2418");
    rule rule_3075;
        ChannelMessage t;
        t <- mod_2411.get(0);
        mod_2410.put(1, t);
    endrule
    rule rule_3076;
        ChannelMessage t;
        t <- mod_2380.get(0);
        mod_2381.put(0, t);
    endrule
    rule rule_3077;
        ChannelMessage t;
        t <- mod_2401.get(0);
        mod_2400.put(0, t);
    endrule
    rule rule_3078;
        ChannelMessage t;
        t <- mod_2412.get(1);
        mod_2387.put(1, t);
    endrule
    rule rule_3079;
        ChannelMessage t;
        t <- mod_2414.get(0);
        mod_2412.put(0, t);
    endrule
    rule rule_3080;
        ChannelMessage t;
        t <- mod_2390.get(0);
        mod_2402.put(0, t);
    endrule
    rule rule_3081;
        ChannelMessage t;
        t <- mod_2393.get(1);
        mod_2394.put(0, t);
    endrule
    rule rule_3082;
        ChannelMessage t;
        t <- mod_2409.get(0);
        mod_2408.put(0, t);
    endrule
    rule rule_3083;
        ChannelMessage t;
        t <- mod_2406.get(1);
        mod_2405.put(1, t);
    endrule
    rule rule_3084;
        ChannelMessage t;
        t <- mod_2385.get(1);
        mod_2386.put(0, t);
    endrule
    rule rule_3085;
        ChannelMessage t;
        t <- mod_2381.get(0);
        mod_2382.put(0, t);
    endrule
    rule rule_3086;
        ChannelMessage t;
        t <- mod_2402.get(0);
        mod_2390.put(1, t);
    endrule
    rule rule_3087;
        ChannelMessage t;
        t <- mod_2394.get(0);
        mod_2396.put(0, t);
    endrule
    rule rule_3088;
        ChannelMessage t;
        t <- mod_2403.get(0);
        mod_2389.put(1, t);
    endrule
    rule rule_3089;
        ChannelMessage t;
        t <- mod_2418.get(0);
        mod_2418.put(1, t);
    endrule
    rule rule_3090;
        ChannelMessage t;
        t <- mod_2396.get(1);
        mod_2394.put(1, t);
    endrule
    rule rule_3091;
        ChannelMessage t;
        t <- mod_2405.get(0);
        mod_2404.put(0, t);
    endrule
    rule rule_3092;
        ChannelMessage t;
        t <- mod_2413.get(0);
        mod_2412.put(1, t);
    endrule
    rule rule_3093;
        ChannelMessage t;
        t <- mod_2404.get(0);
        mod_2403.put(0, t);
    endrule
    rule rule_3094;
        ChannelMessage t;
        t <- mod_2398.get(0);
        mod_2399.put(0, t);
    endrule
    rule rule_3095;
        ChannelMessage t;
        t <- mod_2384.get(1);
        mod_2385.put(0, t);
    endrule
    rule rule_3096;
        ChannelMessage t;
        t <- mod_2389.get(0);
        mod_2390.put(0, t);
    endrule
    rule rule_3097;
        ChannelMessage t;
        t <- mod_2410.get(1);
        mod_2405.put(0, t);
    endrule
    rule rule_3098;
        ChannelMessage t;
        t <- mod_2410.get(0);
        mod_2411.put(0, t);
    endrule
    rule rule_3099;
        ChannelMessage t;
        t <- mod_2385.get(0);
        mod_2410.put(0, t);
    endrule
    rule rule_3100;
        ChannelMessage t;
        t <- mod_2396.get(0);
        mod_2396.put(1, t);
    endrule
    rule rule_3101;
        ChannelMessage t;
        t <- mod_2416.get(0);
        mod_2386.put(1, t);
    endrule
    rule rule_3102;
        ChannelMessage t;
        t <- mod_2386.get(1);
        mod_2387.put(0, t);
    endrule
    rule rule_3103;
        ChannelMessage t;
        t <- mod_2400.get(0);
        mod_2398.put(0, t);
    endrule
    rule rule_3104;
        ChannelMessage t;
        t <- mod_2397.get(1);
        mod_2393.put(1, t);
    endrule
    rule rule_3105;
        ChannelMessage t;
        t <- mod_2415.get(0);
        mod_2414.put(0, t);
    endrule
    rule rule_3106;
        ChannelMessage t;
        t <- mod_2412.get(0);
        mod_2413.put(0, t);
    endrule
    rule rule_3107;
        ChannelMessage t;
        t <- mod_2384.get(0);
        mod_2417.put(0, t);
    endrule
    rule rule_3108;
        ChannelMessage t;
        t <- mod_2387.get(0);
        mod_2388.put(0, t);
    endrule
    rule rule_3109;
        ChannelMessage t;
        t <- mod_2393.get(0);
        mod_2397.put(0, t);
    endrule
    rule rule_3110;
        ChannelMessage t;
        t <- mod_2379.get(0);
        mod_2380.put(0, t);
    endrule
    rule rule_3111;
        ChannelMessage t;
        t <- mod_2417.get(0);
        mod_2384.put(1, t);
    endrule
    rule rule_3112;
        ChannelMessage t;
        t <- mod_2392.get(0);
        mod_2393.put(0, t);
    endrule
    rule rule_3113;
        ChannelMessage t;
        t <- mod_2397.get(0);
        mod_2397.put(1, t);
    endrule
    rule rule_3114;
        ChannelMessage t;
        t <- mod_2388.get(0);
        mod_2389.put(0, t);
    endrule
    rule rule_3115;
        ChannelMessage t;
        t <- mod_2383.get(3);
        mod_2384.put(0, t);
    endrule
    rule rule_3116;
        ChannelMessage t;
        t <- mod_2391.get(0);
        mod_2392.put(0, t);
    endrule
    rule rule_3117;
        ChannelMessage t;
        t <- mod_2382.get(0);
        mod_2418.put(0, t);
    endrule
    rule rule_3118;
        ChannelMessage t;
        t <- mod_2394.get(1);
        mod_2395.put(1, t);
    endrule
    rule rule_3119;
        ChannelMessage t;
        t <- mod_2418.get(1);
        mod_2382.put(1, t);
    endrule
    rule rule_3120;
        ChannelMessage t;
        t <- mod_2407.get(0);
        mod_2406.put(1, t);
    endrule
    rule rule_3121;
        ChannelMessage t;
        t <- mod_2390.get(1);
        mod_2391.put(0, t);
    endrule
    rule rule_3122;
        ChannelMessage t;
        t <- mod_2408.get(0);
        mod_2406.put(0, t);
    endrule
    rule rule_3123;
        ChannelMessage t;
        t <- mod_2399.get(0);
        mod_2398.put(1, t);
    endrule
    rule rule_3124;
        ChannelMessage t;
        t <- mod_2386.get(0);
        mod_2416.put(0, t);
    endrule
    rule rule_3125;
        ChannelMessage t;
        t <- mod_2398.get(1);
        mod_2391.put(1, t);
    endrule
    rule rule_3126;
        ChannelMessage t;
        t <- mod_2406.get(0);
        mod_2407.put(0, t);
    endrule
    rule rule_3127;
        ChannelMessage t;
        t <- mod_2382.get(1);
        mod_2383.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2379.put(0, t);
        end
        if (i == 1) begin
            mod_2395.put(0, t);
        end
        if (i == 2) begin
            mod_2401.put(0, t);
        end
        if (i == 3) begin
            mod_2409.put(0, t);
        end
        if (i == 4) begin
            mod_2415.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_2383.get(0);
        end
        if (i == 3) begin
            t <- mod_2383.get(1);
        end
        if (i == 0) begin
            t <- mod_2383.get(2);
        end
        if (i == 2) begin
            t <- mod_2395.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6093 (Operation_IFC);
    Operation_IFC mod_2420_inner <- mkReshape(2, 64);
    Operation_IFC mod_2420 <- mkDebugOperation(mod_2420_inner, "mod_2420");
    Operation_IFC mod_2421_inner <- mkFlatten(1);
    Operation_IFC mod_2421 <- mkDebugOperation(mod_2421_inner, "mod_2421");
    Operation_IFC mod_2422_inner <- mkFlatten(2);
    Operation_IFC mod_2422 <- mkDebugOperation(mod_2422_inner, "mod_2422");
    Operation_IFC mod_2423_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2423 <- mkDebugOperation(mod_2423_inner, "mod_2423");
    Broadcast_IFC#(4) mod_2424_inner <- mkBroadcast(4);
    Operation_IFC mod_2424 <- mkDebugOperation(mod_2424_inner.op, "mod_2424");
    PMU_IFC mod_2425_bufferize <- mkPMU(2);
    Operation_IFC mod_2425_inner = mod_2425_bufferize.operation;
    Operation_IFC mod_2425 <- mkDebugOperation(mod_2425_inner, "mod_2425");
    Broadcast_IFC#(2) mod_2426_inner <- mkBroadcast(2);
    Operation_IFC mod_2426 <- mkDebugOperation(mod_2426_inner.op, "mod_2426");
    PMU_IFC mod_2427_bufferize <- mkPMU(1);
    Operation_IFC mod_2427_inner = mod_2427_bufferize.operation;
    Operation_IFC mod_2427 <- mkDebugOperation(mod_2427_inner, "mod_2427");
    Operation_IFC mod_2428_inner <- mkBinaryMap(1097, matmul_t_tile);
    Operation_IFC mod_2428 <- mkDebugOperation(mod_2428_inner, "mod_2428");
    Operation_IFC mod_2429_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2429 <- mkDebugOperation(mod_2429_inner, "mod_2429");
    Operation_IFC mod_2430_inner <- mkBinaryMap(1865, mul_tile);
    Operation_IFC mod_2430 <- mkDebugOperation(mod_2430_inner, "mod_2430");
    PMU_IFC mod_2431_bufferize <- mkPMU(1);
    Operation_IFC mod_2431_inner = mod_2431_bufferize.operation;
    Operation_IFC mod_2431 <- mkDebugOperation(mod_2431_inner, "mod_2431");
    Operation_IFC mod_2432_inner <- mkBinaryMap(2445, matmul_t_tile);
    Operation_IFC mod_2432 <- mkDebugOperation(mod_2432_inner, "mod_2432");
    Operation_IFC mod_2433_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2433 <- mkDebugOperation(mod_2433_inner, "mod_2433");
    Operation_IFC mod_2434_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2434 <- mkDebugOperation(mod_2434_inner, "mod_2434");
    Operation_IFC mod_2435_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2435 <- mkDebugOperation(mod_2435_inner, "mod_2435");
    Operation_IFC mod_2436_inner <- mkBinaryMap(2764, mul_tile);
    Operation_IFC mod_2436 <- mkDebugOperation(mod_2436_inner, "mod_2436");
    PMU_IFC mod_2437_bufferize <- mkPMU(1);
    Operation_IFC mod_2437_inner = mod_2437_bufferize.operation;
    Operation_IFC mod_2437 <- mkDebugOperation(mod_2437_inner, "mod_2437");
    PMU_IFC mod_2438_bufferize <- mkPMU(2);
    Operation_IFC mod_2438_inner = mod_2438_bufferize.operation;
    Operation_IFC mod_2438 <- mkDebugOperation(mod_2438_inner, "mod_2438");
    PMU_IFC mod_2439_bufferize <- mkPMU(2);
    Operation_IFC mod_2439_inner = mod_2439_bufferize.operation;
    Operation_IFC mod_2439 <- mkDebugOperation(mod_2439_inner, "mod_2439");
    Operation_IFC mod_2440_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2440 <- mkDebugOperation(mod_2440_inner, "mod_2440");
    Operation_IFC mod_2441_inner <- mkFlatten(1);
    Operation_IFC mod_2441 <- mkDebugOperation(mod_2441_inner, "mod_2441");
    Operation_IFC mod_2442_inner <- mkFlatten(0);
    Operation_IFC mod_2442 <- mkDebugOperation(mod_2442_inner, "mod_2442");
    Operation_IFC mod_2443_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2443 <- mkDebugOperation(mod_2443_inner, "mod_2443");
    Operation_IFC mod_2444_inner <- mkUnaryMap(1737, silu_tile);
    Operation_IFC mod_2444 <- mkDebugOperation(mod_2444_inner, "mod_2444");
    Operation_IFC mod_2445_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2445 <- mkDebugOperation(mod_2445_inner, "mod_2445");
    Operation_IFC mod_2446_inner <- mkBinaryMap(1609, matmul_t_tile);
    Operation_IFC mod_2446 <- mkDebugOperation(mod_2446_inner, "mod_2446");
    PMU_IFC mod_2447_bufferize <- mkPMU(2);
    Operation_IFC mod_2447_inner = mod_2447_bufferize.operation;
    Operation_IFC mod_2447 <- mkDebugOperation(mod_2447_inner, "mod_2447");
    Operation_IFC mod_2448_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2448 <- mkDebugOperation(mod_2448_inner, "mod_2448");
    Operation_IFC mod_2449_inner <- mkFlatten(1);
    Operation_IFC mod_2449 <- mkDebugOperation(mod_2449_inner, "mod_2449");
    Operation_IFC mod_2450_inner <- mkFlatten(0);
    Operation_IFC mod_2450 <- mkDebugOperation(mod_2450_inner, "mod_2450");
    PMU_IFC mod_2451_bufferize <- mkPMU(1);
    Operation_IFC mod_2451_inner = mod_2451_bufferize.operation;
    Operation_IFC mod_2451 <- mkDebugOperation(mod_2451_inner, "mod_2451");
    Operation_IFC mod_2452_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2452 <- mkDebugOperation(mod_2452_inner, "mod_2452");
    PMU_IFC mod_2453_bufferize <- mkPMU(2);
    Operation_IFC mod_2453_inner = mod_2453_bufferize.operation;
    Operation_IFC mod_2453 <- mkDebugOperation(mod_2453_inner, "mod_2453");
    Operation_IFC mod_2454_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2454 <- mkDebugOperation(mod_2454_inner, "mod_2454");
    Operation_IFC mod_2455_inner <- mkFlatten(1);
    Operation_IFC mod_2455 <- mkDebugOperation(mod_2455_inner, "mod_2455");
    Operation_IFC mod_2456_inner <- mkFlatten(0);
    Operation_IFC mod_2456 <- mkDebugOperation(mod_2456_inner, "mod_2456");
    Operation_IFC mod_2457_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2457 <- mkDebugOperation(mod_2457_inner, "mod_2457");
    Operation_IFC mod_2458_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2458 <- mkDebugOperation(mod_2458_inner, "mod_2458");
    PMU_IFC mod_2459_bufferize <- mkPMU(2);
    Operation_IFC mod_2459_inner = mod_2459_bufferize.operation;
    Operation_IFC mod_2459 <- mkDebugOperation(mod_2459_inner, "mod_2459");
    rule rule_3128;
        ChannelMessage t;
        t <- mod_2447.get(1);
        mod_2446.put(1, t);
    endrule
    rule rule_3129;
        ChannelMessage t;
        t <- mod_2449.get(0);
        mod_2447.put(0, t);
    endrule
    rule rule_3130;
        ChannelMessage t;
        t <- mod_2431.get(0);
        mod_2443.put(0, t);
    endrule
    rule rule_3131;
        ChannelMessage t;
        t <- mod_2447.get(0);
        mod_2448.put(0, t);
    endrule
    rule rule_3132;
        ChannelMessage t;
        t <- mod_2425.get(1);
        mod_2426.put(0, t);
    endrule
    rule rule_3133;
        ChannelMessage t;
        t <- mod_2427.get(1);
        mod_2428.put(0, t);
    endrule
    rule rule_3134;
        ChannelMessage t;
        t <- mod_2451.get(0);
        mod_2452.put(0, t);
    endrule
    rule rule_3135;
        ChannelMessage t;
        t <- mod_2434.get(0);
        mod_2438.put(0, t);
    endrule
    rule rule_3136;
        ChannelMessage t;
        t <- mod_2453.get(1);
        mod_2428.put(1, t);
    endrule
    rule rule_3137;
        ChannelMessage t;
        t <- mod_2450.get(0);
        mod_2449.put(0, t);
    endrule
    rule rule_3138;
        ChannelMessage t;
        t <- mod_2433.get(0);
        mod_2434.put(0, t);
    endrule
    rule rule_3139;
        ChannelMessage t;
        t <- mod_2457.get(0);
        mod_2427.put(1, t);
    endrule
    rule rule_3140;
        ChannelMessage t;
        t <- mod_2424.get(3);
        mod_2425.put(0, t);
    endrule
    rule rule_3141;
        ChannelMessage t;
        t <- mod_2446.get(0);
        mod_2445.put(0, t);
    endrule
    rule rule_3142;
        ChannelMessage t;
        t <- mod_2439.get(0);
        mod_2440.put(0, t);
    endrule
    rule rule_3143;
        ChannelMessage t;
        t <- mod_2456.get(0);
        mod_2455.put(0, t);
    endrule
    rule rule_3144;
        ChannelMessage t;
        t <- mod_2458.get(0);
        mod_2425.put(1, t);
    endrule
    rule rule_3145;
        ChannelMessage t;
        t <- mod_2427.get(0);
        mod_2457.put(0, t);
    endrule
    rule rule_3146;
        ChannelMessage t;
        t <- mod_2420.get(0);
        mod_2421.put(0, t);
    endrule
    rule rule_3147;
        ChannelMessage t;
        t <- mod_2422.get(0);
        mod_2423.put(0, t);
    endrule
    rule rule_3148;
        ChannelMessage t;
        t <- mod_2437.get(1);
        mod_2435.put(1, t);
    endrule
    rule rule_3149;
        ChannelMessage t;
        t <- mod_2435.get(0);
        mod_2437.put(0, t);
    endrule
    rule rule_3150;
        ChannelMessage t;
        t <- mod_2426.get(0);
        mod_2451.put(0, t);
    endrule
    rule rule_3151;
        ChannelMessage t;
        t <- mod_2435.get(1);
        mod_2436.put(1, t);
    endrule
    rule rule_3152;
        ChannelMessage t;
        t <- mod_2438.get(1);
        mod_2434.put(1, t);
    endrule
    rule rule_3153;
        ChannelMessage t;
        t <- mod_2440.get(0);
        mod_2439.put(1, t);
    endrule
    rule rule_3154;
        ChannelMessage t;
        t <- mod_2448.get(0);
        mod_2447.put(1, t);
    endrule
    rule rule_3155;
        ChannelMessage t;
        t <- mod_2441.get(0);
        mod_2439.put(0, t);
    endrule
    rule rule_3156;
        ChannelMessage t;
        t <- mod_2434.get(1);
        mod_2435.put(0, t);
    endrule
    rule rule_3157;
        ChannelMessage t;
        t <- mod_2437.get(0);
        mod_2437.put(1, t);
    endrule
    rule rule_3158;
        ChannelMessage t;
        t <- mod_2421.get(0);
        mod_2422.put(0, t);
    endrule
    rule rule_3159;
        ChannelMessage t;
        t <- mod_2455.get(0);
        mod_2453.put(0, t);
    endrule
    rule rule_3160;
        ChannelMessage t;
        t <- mod_2438.get(0);
        mod_2438.put(1, t);
    endrule
    rule rule_3161;
        ChannelMessage t;
        t <- mod_2430.get(0);
        mod_2431.put(0, t);
    endrule
    rule rule_3162;
        ChannelMessage t;
        t <- mod_2432.get(0);
        mod_2433.put(0, t);
    endrule
    rule rule_3163;
        ChannelMessage t;
        t <- mod_2444.get(0);
        mod_2430.put(1, t);
    endrule
    rule rule_3164;
        ChannelMessage t;
        t <- mod_2428.get(0);
        mod_2429.put(0, t);
    endrule
    rule rule_3165;
        ChannelMessage t;
        t <- mod_2439.get(1);
        mod_2432.put(1, t);
    endrule
    rule rule_3166;
        ChannelMessage t;
        t <- mod_2442.get(0);
        mod_2441.put(0, t);
    endrule
    rule rule_3167;
        ChannelMessage t;
        t <- mod_2423.get(1);
        mod_2424.put(0, t);
    endrule
    rule rule_3168;
        ChannelMessage t;
        t <- mod_2429.get(0);
        mod_2430.put(0, t);
    endrule
    rule rule_3169;
        ChannelMessage t;
        t <- mod_2454.get(0);
        mod_2453.put(1, t);
    endrule
    rule rule_3170;
        ChannelMessage t;
        t <- mod_2459.get(0);
        mod_2459.put(1, t);
    endrule
    rule rule_3171;
        ChannelMessage t;
        t <- mod_2453.get(0);
        mod_2454.put(0, t);
    endrule
    rule rule_3172;
        ChannelMessage t;
        t <- mod_2443.get(0);
        mod_2431.put(1, t);
    endrule
    rule rule_3173;
        ChannelMessage t;
        t <- mod_2452.get(0);
        mod_2451.put(1, t);
    endrule
    rule rule_3174;
        ChannelMessage t;
        t <- mod_2451.get(1);
        mod_2446.put(0, t);
    endrule
    rule rule_3175;
        ChannelMessage t;
        t <- mod_2431.get(1);
        mod_2432.put(0, t);
    endrule
    rule rule_3176;
        ChannelMessage t;
        t <- mod_2445.get(0);
        mod_2444.put(0, t);
    endrule
    rule rule_3177;
        ChannelMessage t;
        t <- mod_2459.get(1);
        mod_2423.put(1, t);
    endrule
    rule rule_3178;
        ChannelMessage t;
        t <- mod_2423.get(0);
        mod_2459.put(0, t);
    endrule
    rule rule_3179;
        ChannelMessage t;
        t <- mod_2425.get(0);
        mod_2458.put(0, t);
    endrule
    rule rule_3180;
        ChannelMessage t;
        t <- mod_2426.get(1);
        mod_2427.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2420.put(0, t);
        end
        if (i == 1) begin
            mod_2436.put(0, t);
        end
        if (i == 2) begin
            mod_2442.put(0, t);
        end
        if (i == 3) begin
            mod_2450.put(0, t);
        end
        if (i == 4) begin
            mod_2456.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 2) begin
            t <- mod_2424.get(0);
        end
        if (i == 1) begin
            t <- mod_2424.get(1);
        end
        if (i == 3) begin
            t <- mod_2424.get(2);
        end
        if (i == 0) begin
            t <- mod_2436.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6094 (Operation_IFC);
    Operation_IFC mod_2461_inner <- mkReshape(2, 64);
    Operation_IFC mod_2461 <- mkDebugOperation(mod_2461_inner, "mod_2461");
    Operation_IFC mod_2462_inner <- mkFlatten(1);
    Operation_IFC mod_2462 <- mkDebugOperation(mod_2462_inner, "mod_2462");
    Operation_IFC mod_2463_inner <- mkFlatten(2);
    Operation_IFC mod_2463 <- mkDebugOperation(mod_2463_inner, "mod_2463");
    Operation_IFC mod_2464_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2464 <- mkDebugOperation(mod_2464_inner, "mod_2464");
    Broadcast_IFC#(4) mod_2465_inner <- mkBroadcast(4);
    Operation_IFC mod_2465 <- mkDebugOperation(mod_2465_inner.op, "mod_2465");
    PMU_IFC mod_2466_bufferize <- mkPMU(2);
    Operation_IFC mod_2466_inner = mod_2466_bufferize.operation;
    Operation_IFC mod_2466 <- mkDebugOperation(mod_2466_inner, "mod_2466");
    Broadcast_IFC#(2) mod_2467_inner <- mkBroadcast(2);
    Operation_IFC mod_2467 <- mkDebugOperation(mod_2467_inner.op, "mod_2467");
    PMU_IFC mod_2468_bufferize <- mkPMU(1);
    Operation_IFC mod_2468_inner = mod_2468_bufferize.operation;
    Operation_IFC mod_2468 <- mkDebugOperation(mod_2468_inner, "mod_2468");
    Operation_IFC mod_2469_inner <- mkBinaryMap(1096, matmul_t_tile);
    Operation_IFC mod_2469 <- mkDebugOperation(mod_2469_inner, "mod_2469");
    Operation_IFC mod_2470_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2470 <- mkDebugOperation(mod_2470_inner, "mod_2470");
    Operation_IFC mod_2471_inner <- mkBinaryMap(1864, mul_tile);
    Operation_IFC mod_2471 <- mkDebugOperation(mod_2471_inner, "mod_2471");
    PMU_IFC mod_2472_bufferize <- mkPMU(1);
    Operation_IFC mod_2472_inner = mod_2472_bufferize.operation;
    Operation_IFC mod_2472 <- mkDebugOperation(mod_2472_inner, "mod_2472");
    Operation_IFC mod_2473_inner <- mkBinaryMap(2443, matmul_t_tile);
    Operation_IFC mod_2473 <- mkDebugOperation(mod_2473_inner, "mod_2473");
    Operation_IFC mod_2474_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2474 <- mkDebugOperation(mod_2474_inner, "mod_2474");
    Operation_IFC mod_2475_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2475 <- mkDebugOperation(mod_2475_inner, "mod_2475");
    Operation_IFC mod_2476_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2476 <- mkDebugOperation(mod_2476_inner, "mod_2476");
    Operation_IFC mod_2477_inner <- mkBinaryMap(2763, mul_tile);
    Operation_IFC mod_2477 <- mkDebugOperation(mod_2477_inner, "mod_2477");
    PMU_IFC mod_2478_bufferize <- mkPMU(1);
    Operation_IFC mod_2478_inner = mod_2478_bufferize.operation;
    Operation_IFC mod_2478 <- mkDebugOperation(mod_2478_inner, "mod_2478");
    PMU_IFC mod_2479_bufferize <- mkPMU(2);
    Operation_IFC mod_2479_inner = mod_2479_bufferize.operation;
    Operation_IFC mod_2479 <- mkDebugOperation(mod_2479_inner, "mod_2479");
    PMU_IFC mod_2480_bufferize <- mkPMU(2);
    Operation_IFC mod_2480_inner = mod_2480_bufferize.operation;
    Operation_IFC mod_2480 <- mkDebugOperation(mod_2480_inner, "mod_2480");
    Operation_IFC mod_2481_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2481 <- mkDebugOperation(mod_2481_inner, "mod_2481");
    Operation_IFC mod_2482_inner <- mkFlatten(1);
    Operation_IFC mod_2482 <- mkDebugOperation(mod_2482_inner, "mod_2482");
    Operation_IFC mod_2483_inner <- mkFlatten(0);
    Operation_IFC mod_2483 <- mkDebugOperation(mod_2483_inner, "mod_2483");
    Operation_IFC mod_2484_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2484 <- mkDebugOperation(mod_2484_inner, "mod_2484");
    Operation_IFC mod_2485_inner <- mkUnaryMap(1736, silu_tile);
    Operation_IFC mod_2485 <- mkDebugOperation(mod_2485_inner, "mod_2485");
    Operation_IFC mod_2486_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2486 <- mkDebugOperation(mod_2486_inner, "mod_2486");
    Operation_IFC mod_2487_inner <- mkBinaryMap(1608, matmul_t_tile);
    Operation_IFC mod_2487 <- mkDebugOperation(mod_2487_inner, "mod_2487");
    PMU_IFC mod_2488_bufferize <- mkPMU(2);
    Operation_IFC mod_2488_inner = mod_2488_bufferize.operation;
    Operation_IFC mod_2488 <- mkDebugOperation(mod_2488_inner, "mod_2488");
    Operation_IFC mod_2489_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2489 <- mkDebugOperation(mod_2489_inner, "mod_2489");
    Operation_IFC mod_2490_inner <- mkFlatten(1);
    Operation_IFC mod_2490 <- mkDebugOperation(mod_2490_inner, "mod_2490");
    Operation_IFC mod_2491_inner <- mkFlatten(0);
    Operation_IFC mod_2491 <- mkDebugOperation(mod_2491_inner, "mod_2491");
    PMU_IFC mod_2492_bufferize <- mkPMU(1);
    Operation_IFC mod_2492_inner = mod_2492_bufferize.operation;
    Operation_IFC mod_2492 <- mkDebugOperation(mod_2492_inner, "mod_2492");
    Operation_IFC mod_2493_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2493 <- mkDebugOperation(mod_2493_inner, "mod_2493");
    PMU_IFC mod_2494_bufferize <- mkPMU(2);
    Operation_IFC mod_2494_inner = mod_2494_bufferize.operation;
    Operation_IFC mod_2494 <- mkDebugOperation(mod_2494_inner, "mod_2494");
    Operation_IFC mod_2495_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2495 <- mkDebugOperation(mod_2495_inner, "mod_2495");
    Operation_IFC mod_2496_inner <- mkFlatten(1);
    Operation_IFC mod_2496 <- mkDebugOperation(mod_2496_inner, "mod_2496");
    Operation_IFC mod_2497_inner <- mkFlatten(0);
    Operation_IFC mod_2497 <- mkDebugOperation(mod_2497_inner, "mod_2497");
    Operation_IFC mod_2498_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2498 <- mkDebugOperation(mod_2498_inner, "mod_2498");
    Operation_IFC mod_2499_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2499 <- mkDebugOperation(mod_2499_inner, "mod_2499");
    PMU_IFC mod_2500_bufferize <- mkPMU(2);
    Operation_IFC mod_2500_inner = mod_2500_bufferize.operation;
    Operation_IFC mod_2500 <- mkDebugOperation(mod_2500_inner, "mod_2500");
    rule rule_3181;
        ChannelMessage t;
        t <- mod_2474.get(0);
        mod_2475.put(0, t);
    endrule
    rule rule_3182;
        ChannelMessage t;
        t <- mod_2482.get(0);
        mod_2480.put(0, t);
    endrule
    rule rule_3183;
        ChannelMessage t;
        t <- mod_2489.get(0);
        mod_2488.put(1, t);
    endrule
    rule rule_3184;
        ChannelMessage t;
        t <- mod_2491.get(0);
        mod_2490.put(0, t);
    endrule
    rule rule_3185;
        ChannelMessage t;
        t <- mod_2479.get(0);
        mod_2479.put(1, t);
    endrule
    rule rule_3186;
        ChannelMessage t;
        t <- mod_2476.get(0);
        mod_2478.put(0, t);
    endrule
    rule rule_3187;
        ChannelMessage t;
        t <- mod_2490.get(0);
        mod_2488.put(0, t);
    endrule
    rule rule_3188;
        ChannelMessage t;
        t <- mod_2492.get(1);
        mod_2487.put(0, t);
    endrule
    rule rule_3189;
        ChannelMessage t;
        t <- mod_2486.get(0);
        mod_2485.put(0, t);
    endrule
    rule rule_3190;
        ChannelMessage t;
        t <- mod_2468.get(1);
        mod_2469.put(0, t);
    endrule
    rule rule_3191;
        ChannelMessage t;
        t <- mod_2500.get(0);
        mod_2500.put(1, t);
    endrule
    rule rule_3192;
        ChannelMessage t;
        t <- mod_2488.get(0);
        mod_2489.put(0, t);
    endrule
    rule rule_3193;
        ChannelMessage t;
        t <- mod_2480.get(1);
        mod_2473.put(1, t);
    endrule
    rule rule_3194;
        ChannelMessage t;
        t <- mod_2494.get(1);
        mod_2469.put(1, t);
    endrule
    rule rule_3195;
        ChannelMessage t;
        t <- mod_2498.get(0);
        mod_2468.put(1, t);
    endrule
    rule rule_3196;
        ChannelMessage t;
        t <- mod_2475.get(0);
        mod_2479.put(0, t);
    endrule
    rule rule_3197;
        ChannelMessage t;
        t <- mod_2467.get(1);
        mod_2468.put(0, t);
    endrule
    rule rule_3198;
        ChannelMessage t;
        t <- mod_2468.get(0);
        mod_2498.put(0, t);
    endrule
    rule rule_3199;
        ChannelMessage t;
        t <- mod_2483.get(0);
        mod_2482.put(0, t);
    endrule
    rule rule_3200;
        ChannelMessage t;
        t <- mod_2470.get(0);
        mod_2471.put(0, t);
    endrule
    rule rule_3201;
        ChannelMessage t;
        t <- mod_2461.get(0);
        mod_2462.put(0, t);
    endrule
    rule rule_3202;
        ChannelMessage t;
        t <- mod_2464.get(1);
        mod_2465.put(0, t);
    endrule
    rule rule_3203;
        ChannelMessage t;
        t <- mod_2469.get(0);
        mod_2470.put(0, t);
    endrule
    rule rule_3204;
        ChannelMessage t;
        t <- mod_2476.get(1);
        mod_2477.put(1, t);
    endrule
    rule rule_3205;
        ChannelMessage t;
        t <- mod_2496.get(0);
        mod_2494.put(0, t);
    endrule
    rule rule_3206;
        ChannelMessage t;
        t <- mod_2471.get(0);
        mod_2472.put(0, t);
    endrule
    rule rule_3207;
        ChannelMessage t;
        t <- mod_2484.get(0);
        mod_2472.put(1, t);
    endrule
    rule rule_3208;
        ChannelMessage t;
        t <- mod_2472.get(1);
        mod_2473.put(0, t);
    endrule
    rule rule_3209;
        ChannelMessage t;
        t <- mod_2500.get(1);
        mod_2464.put(1, t);
    endrule
    rule rule_3210;
        ChannelMessage t;
        t <- mod_2493.get(0);
        mod_2492.put(1, t);
    endrule
    rule rule_3211;
        ChannelMessage t;
        t <- mod_2466.get(0);
        mod_2499.put(0, t);
    endrule
    rule rule_3212;
        ChannelMessage t;
        t <- mod_2478.get(0);
        mod_2478.put(1, t);
    endrule
    rule rule_3213;
        ChannelMessage t;
        t <- mod_2464.get(0);
        mod_2500.put(0, t);
    endrule
    rule rule_3214;
        ChannelMessage t;
        t <- mod_2467.get(0);
        mod_2492.put(0, t);
    endrule
    rule rule_3215;
        ChannelMessage t;
        t <- mod_2475.get(1);
        mod_2476.put(0, t);
    endrule
    rule rule_3216;
        ChannelMessage t;
        t <- mod_2494.get(0);
        mod_2495.put(0, t);
    endrule
    rule rule_3217;
        ChannelMessage t;
        t <- mod_2492.get(0);
        mod_2493.put(0, t);
    endrule
    rule rule_3218;
        ChannelMessage t;
        t <- mod_2488.get(1);
        mod_2487.put(1, t);
    endrule
    rule rule_3219;
        ChannelMessage t;
        t <- mod_2495.get(0);
        mod_2494.put(1, t);
    endrule
    rule rule_3220;
        ChannelMessage t;
        t <- mod_2479.get(1);
        mod_2475.put(1, t);
    endrule
    rule rule_3221;
        ChannelMessage t;
        t <- mod_2465.get(3);
        mod_2466.put(0, t);
    endrule
    rule rule_3222;
        ChannelMessage t;
        t <- mod_2478.get(1);
        mod_2476.put(1, t);
    endrule
    rule rule_3223;
        ChannelMessage t;
        t <- mod_2485.get(0);
        mod_2471.put(1, t);
    endrule
    rule rule_3224;
        ChannelMessage t;
        t <- mod_2462.get(0);
        mod_2463.put(0, t);
    endrule
    rule rule_3225;
        ChannelMessage t;
        t <- mod_2480.get(0);
        mod_2481.put(0, t);
    endrule
    rule rule_3226;
        ChannelMessage t;
        t <- mod_2472.get(0);
        mod_2484.put(0, t);
    endrule
    rule rule_3227;
        ChannelMessage t;
        t <- mod_2481.get(0);
        mod_2480.put(1, t);
    endrule
    rule rule_3228;
        ChannelMessage t;
        t <- mod_2473.get(0);
        mod_2474.put(0, t);
    endrule
    rule rule_3229;
        ChannelMessage t;
        t <- mod_2463.get(0);
        mod_2464.put(0, t);
    endrule
    rule rule_3230;
        ChannelMessage t;
        t <- mod_2499.get(0);
        mod_2466.put(1, t);
    endrule
    rule rule_3231;
        ChannelMessage t;
        t <- mod_2466.get(1);
        mod_2467.put(0, t);
    endrule
    rule rule_3232;
        ChannelMessage t;
        t <- mod_2487.get(0);
        mod_2486.put(0, t);
    endrule
    rule rule_3233;
        ChannelMessage t;
        t <- mod_2497.get(0);
        mod_2496.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2461.put(0, t);
        end
        if (i == 1) begin
            mod_2477.put(0, t);
        end
        if (i == 2) begin
            mod_2483.put(0, t);
        end
        if (i == 3) begin
            mod_2491.put(0, t);
        end
        if (i == 4) begin
            mod_2497.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_2465.get(0);
        end
        if (i == 2) begin
            t <- mod_2465.get(1);
        end
        if (i == 3) begin
            t <- mod_2465.get(2);
        end
        if (i == 0) begin
            t <- mod_2477.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6095 (Operation_IFC);
    Operation_IFC mod_2502_inner <- mkReshape(2, 64);
    Operation_IFC mod_2502 <- mkDebugOperation(mod_2502_inner, "mod_2502");
    Operation_IFC mod_2503_inner <- mkFlatten(1);
    Operation_IFC mod_2503 <- mkDebugOperation(mod_2503_inner, "mod_2503");
    Operation_IFC mod_2504_inner <- mkFlatten(2);
    Operation_IFC mod_2504 <- mkDebugOperation(mod_2504_inner, "mod_2504");
    Operation_IFC mod_2505_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2505 <- mkDebugOperation(mod_2505_inner, "mod_2505");
    Broadcast_IFC#(4) mod_2506_inner <- mkBroadcast(4);
    Operation_IFC mod_2506 <- mkDebugOperation(mod_2506_inner.op, "mod_2506");
    PMU_IFC mod_2507_bufferize <- mkPMU(2);
    Operation_IFC mod_2507_inner = mod_2507_bufferize.operation;
    Operation_IFC mod_2507 <- mkDebugOperation(mod_2507_inner, "mod_2507");
    Broadcast_IFC#(2) mod_2508_inner <- mkBroadcast(2);
    Operation_IFC mod_2508 <- mkDebugOperation(mod_2508_inner.op, "mod_2508");
    PMU_IFC mod_2509_bufferize <- mkPMU(1);
    Operation_IFC mod_2509_inner = mod_2509_bufferize.operation;
    Operation_IFC mod_2509 <- mkDebugOperation(mod_2509_inner, "mod_2509");
    Operation_IFC mod_2510_inner <- mkBinaryMap(1095, matmul_t_tile);
    Operation_IFC mod_2510 <- mkDebugOperation(mod_2510_inner, "mod_2510");
    Operation_IFC mod_2511_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2511 <- mkDebugOperation(mod_2511_inner, "mod_2511");
    Operation_IFC mod_2512_inner <- mkBinaryMap(1863, mul_tile);
    Operation_IFC mod_2512 <- mkDebugOperation(mod_2512_inner, "mod_2512");
    PMU_IFC mod_2513_bufferize <- mkPMU(1);
    Operation_IFC mod_2513_inner = mod_2513_bufferize.operation;
    Operation_IFC mod_2513 <- mkDebugOperation(mod_2513_inner, "mod_2513");
    Operation_IFC mod_2514_inner <- mkBinaryMap(2441, matmul_t_tile);
    Operation_IFC mod_2514 <- mkDebugOperation(mod_2514_inner, "mod_2514");
    Operation_IFC mod_2515_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2515 <- mkDebugOperation(mod_2515_inner, "mod_2515");
    Operation_IFC mod_2516_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2516 <- mkDebugOperation(mod_2516_inner, "mod_2516");
    Operation_IFC mod_2517_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2517 <- mkDebugOperation(mod_2517_inner, "mod_2517");
    Operation_IFC mod_2518_inner <- mkBinaryMap(2762, mul_tile);
    Operation_IFC mod_2518 <- mkDebugOperation(mod_2518_inner, "mod_2518");
    PMU_IFC mod_2519_bufferize <- mkPMU(1);
    Operation_IFC mod_2519_inner = mod_2519_bufferize.operation;
    Operation_IFC mod_2519 <- mkDebugOperation(mod_2519_inner, "mod_2519");
    PMU_IFC mod_2520_bufferize <- mkPMU(2);
    Operation_IFC mod_2520_inner = mod_2520_bufferize.operation;
    Operation_IFC mod_2520 <- mkDebugOperation(mod_2520_inner, "mod_2520");
    PMU_IFC mod_2521_bufferize <- mkPMU(2);
    Operation_IFC mod_2521_inner = mod_2521_bufferize.operation;
    Operation_IFC mod_2521 <- mkDebugOperation(mod_2521_inner, "mod_2521");
    Operation_IFC mod_2522_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2522 <- mkDebugOperation(mod_2522_inner, "mod_2522");
    Operation_IFC mod_2523_inner <- mkFlatten(1);
    Operation_IFC mod_2523 <- mkDebugOperation(mod_2523_inner, "mod_2523");
    Operation_IFC mod_2524_inner <- mkFlatten(0);
    Operation_IFC mod_2524 <- mkDebugOperation(mod_2524_inner, "mod_2524");
    Operation_IFC mod_2525_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2525 <- mkDebugOperation(mod_2525_inner, "mod_2525");
    Operation_IFC mod_2526_inner <- mkUnaryMap(1735, silu_tile);
    Operation_IFC mod_2526 <- mkDebugOperation(mod_2526_inner, "mod_2526");
    Operation_IFC mod_2527_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2527 <- mkDebugOperation(mod_2527_inner, "mod_2527");
    Operation_IFC mod_2528_inner <- mkBinaryMap(1607, matmul_t_tile);
    Operation_IFC mod_2528 <- mkDebugOperation(mod_2528_inner, "mod_2528");
    PMU_IFC mod_2529_bufferize <- mkPMU(2);
    Operation_IFC mod_2529_inner = mod_2529_bufferize.operation;
    Operation_IFC mod_2529 <- mkDebugOperation(mod_2529_inner, "mod_2529");
    Operation_IFC mod_2530_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2530 <- mkDebugOperation(mod_2530_inner, "mod_2530");
    Operation_IFC mod_2531_inner <- mkFlatten(1);
    Operation_IFC mod_2531 <- mkDebugOperation(mod_2531_inner, "mod_2531");
    Operation_IFC mod_2532_inner <- mkFlatten(0);
    Operation_IFC mod_2532 <- mkDebugOperation(mod_2532_inner, "mod_2532");
    PMU_IFC mod_2533_bufferize <- mkPMU(1);
    Operation_IFC mod_2533_inner = mod_2533_bufferize.operation;
    Operation_IFC mod_2533 <- mkDebugOperation(mod_2533_inner, "mod_2533");
    Operation_IFC mod_2534_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2534 <- mkDebugOperation(mod_2534_inner, "mod_2534");
    PMU_IFC mod_2535_bufferize <- mkPMU(2);
    Operation_IFC mod_2535_inner = mod_2535_bufferize.operation;
    Operation_IFC mod_2535 <- mkDebugOperation(mod_2535_inner, "mod_2535");
    Operation_IFC mod_2536_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2536 <- mkDebugOperation(mod_2536_inner, "mod_2536");
    Operation_IFC mod_2537_inner <- mkFlatten(1);
    Operation_IFC mod_2537 <- mkDebugOperation(mod_2537_inner, "mod_2537");
    Operation_IFC mod_2538_inner <- mkFlatten(0);
    Operation_IFC mod_2538 <- mkDebugOperation(mod_2538_inner, "mod_2538");
    Operation_IFC mod_2539_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2539 <- mkDebugOperation(mod_2539_inner, "mod_2539");
    Operation_IFC mod_2540_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2540 <- mkDebugOperation(mod_2540_inner, "mod_2540");
    PMU_IFC mod_2541_bufferize <- mkPMU(2);
    Operation_IFC mod_2541_inner = mod_2541_bufferize.operation;
    Operation_IFC mod_2541 <- mkDebugOperation(mod_2541_inner, "mod_2541");
    rule rule_3234;
        ChannelMessage t;
        t <- mod_2540.get(0);
        mod_2507.put(1, t);
    endrule
    rule rule_3235;
        ChannelMessage t;
        t <- mod_2517.get(0);
        mod_2519.put(0, t);
    endrule
    rule rule_3236;
        ChannelMessage t;
        t <- mod_2532.get(0);
        mod_2531.put(0, t);
    endrule
    rule rule_3237;
        ChannelMessage t;
        t <- mod_2507.get(0);
        mod_2540.put(0, t);
    endrule
    rule rule_3238;
        ChannelMessage t;
        t <- mod_2528.get(0);
        mod_2527.put(0, t);
    endrule
    rule rule_3239;
        ChannelMessage t;
        t <- mod_2535.get(0);
        mod_2536.put(0, t);
    endrule
    rule rule_3240;
        ChannelMessage t;
        t <- mod_2538.get(0);
        mod_2537.put(0, t);
    endrule
    rule rule_3241;
        ChannelMessage t;
        t <- mod_2533.get(0);
        mod_2534.put(0, t);
    endrule
    rule rule_3242;
        ChannelMessage t;
        t <- mod_2522.get(0);
        mod_2521.put(1, t);
    endrule
    rule rule_3243;
        ChannelMessage t;
        t <- mod_2531.get(0);
        mod_2529.put(0, t);
    endrule
    rule rule_3244;
        ChannelMessage t;
        t <- mod_2502.get(0);
        mod_2503.put(0, t);
    endrule
    rule rule_3245;
        ChannelMessage t;
        t <- mod_2509.get(1);
        mod_2510.put(0, t);
    endrule
    rule rule_3246;
        ChannelMessage t;
        t <- mod_2515.get(0);
        mod_2516.put(0, t);
    endrule
    rule rule_3247;
        ChannelMessage t;
        t <- mod_2526.get(0);
        mod_2512.put(1, t);
    endrule
    rule rule_3248;
        ChannelMessage t;
        t <- mod_2527.get(0);
        mod_2526.put(0, t);
    endrule
    rule rule_3249;
        ChannelMessage t;
        t <- mod_2506.get(3);
        mod_2507.put(0, t);
    endrule
    rule rule_3250;
        ChannelMessage t;
        t <- mod_2505.get(0);
        mod_2541.put(0, t);
    endrule
    rule rule_3251;
        ChannelMessage t;
        t <- mod_2517.get(1);
        mod_2518.put(1, t);
    endrule
    rule rule_3252;
        ChannelMessage t;
        t <- mod_2519.get(0);
        mod_2519.put(1, t);
    endrule
    rule rule_3253;
        ChannelMessage t;
        t <- mod_2533.get(1);
        mod_2528.put(0, t);
    endrule
    rule rule_3254;
        ChannelMessage t;
        t <- mod_2524.get(0);
        mod_2523.put(0, t);
    endrule
    rule rule_3255;
        ChannelMessage t;
        t <- mod_2534.get(0);
        mod_2533.put(1, t);
    endrule
    rule rule_3256;
        ChannelMessage t;
        t <- mod_2541.get(1);
        mod_2505.put(1, t);
    endrule
    rule rule_3257;
        ChannelMessage t;
        t <- mod_2511.get(0);
        mod_2512.put(0, t);
    endrule
    rule rule_3258;
        ChannelMessage t;
        t <- mod_2512.get(0);
        mod_2513.put(0, t);
    endrule
    rule rule_3259;
        ChannelMessage t;
        t <- mod_2505.get(1);
        mod_2506.put(0, t);
    endrule
    rule rule_3260;
        ChannelMessage t;
        t <- mod_2541.get(0);
        mod_2541.put(1, t);
    endrule
    rule rule_3261;
        ChannelMessage t;
        t <- mod_2519.get(1);
        mod_2517.put(1, t);
    endrule
    rule rule_3262;
        ChannelMessage t;
        t <- mod_2520.get(0);
        mod_2520.put(1, t);
    endrule
    rule rule_3263;
        ChannelMessage t;
        t <- mod_2504.get(0);
        mod_2505.put(0, t);
    endrule
    rule rule_3264;
        ChannelMessage t;
        t <- mod_2525.get(0);
        mod_2513.put(1, t);
    endrule
    rule rule_3265;
        ChannelMessage t;
        t <- mod_2507.get(1);
        mod_2508.put(0, t);
    endrule
    rule rule_3266;
        ChannelMessage t;
        t <- mod_2539.get(0);
        mod_2509.put(1, t);
    endrule
    rule rule_3267;
        ChannelMessage t;
        t <- mod_2530.get(0);
        mod_2529.put(1, t);
    endrule
    rule rule_3268;
        ChannelMessage t;
        t <- mod_2509.get(0);
        mod_2539.put(0, t);
    endrule
    rule rule_3269;
        ChannelMessage t;
        t <- mod_2529.get(0);
        mod_2530.put(0, t);
    endrule
    rule rule_3270;
        ChannelMessage t;
        t <- mod_2513.get(0);
        mod_2525.put(0, t);
    endrule
    rule rule_3271;
        ChannelMessage t;
        t <- mod_2521.get(1);
        mod_2514.put(1, t);
    endrule
    rule rule_3272;
        ChannelMessage t;
        t <- mod_2529.get(1);
        mod_2528.put(1, t);
    endrule
    rule rule_3273;
        ChannelMessage t;
        t <- mod_2536.get(0);
        mod_2535.put(1, t);
    endrule
    rule rule_3274;
        ChannelMessage t;
        t <- mod_2508.get(0);
        mod_2533.put(0, t);
    endrule
    rule rule_3275;
        ChannelMessage t;
        t <- mod_2516.get(1);
        mod_2517.put(0, t);
    endrule
    rule rule_3276;
        ChannelMessage t;
        t <- mod_2537.get(0);
        mod_2535.put(0, t);
    endrule
    rule rule_3277;
        ChannelMessage t;
        t <- mod_2516.get(0);
        mod_2520.put(0, t);
    endrule
    rule rule_3278;
        ChannelMessage t;
        t <- mod_2513.get(1);
        mod_2514.put(0, t);
    endrule
    rule rule_3279;
        ChannelMessage t;
        t <- mod_2503.get(0);
        mod_2504.put(0, t);
    endrule
    rule rule_3280;
        ChannelMessage t;
        t <- mod_2520.get(1);
        mod_2516.put(1, t);
    endrule
    rule rule_3281;
        ChannelMessage t;
        t <- mod_2514.get(0);
        mod_2515.put(0, t);
    endrule
    rule rule_3282;
        ChannelMessage t;
        t <- mod_2510.get(0);
        mod_2511.put(0, t);
    endrule
    rule rule_3283;
        ChannelMessage t;
        t <- mod_2508.get(1);
        mod_2509.put(0, t);
    endrule
    rule rule_3284;
        ChannelMessage t;
        t <- mod_2523.get(0);
        mod_2521.put(0, t);
    endrule
    rule rule_3285;
        ChannelMessage t;
        t <- mod_2521.get(0);
        mod_2522.put(0, t);
    endrule
    rule rule_3286;
        ChannelMessage t;
        t <- mod_2535.get(1);
        mod_2510.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2502.put(0, t);
        end
        if (i == 1) begin
            mod_2518.put(0, t);
        end
        if (i == 2) begin
            mod_2524.put(0, t);
        end
        if (i == 3) begin
            mod_2532.put(0, t);
        end
        if (i == 4) begin
            mod_2538.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 2) begin
            t <- mod_2506.get(0);
        end
        if (i == 1) begin
            t <- mod_2506.get(1);
        end
        if (i == 0) begin
            t <- mod_2506.get(2);
        end
        if (i == 3) begin
            t <- mod_2518.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6096 (Operation_IFC);
    Operation_IFC mod_2543_inner <- mkReshape(2, 64);
    Operation_IFC mod_2543 <- mkDebugOperation(mod_2543_inner, "mod_2543");
    Operation_IFC mod_2544_inner <- mkFlatten(1);
    Operation_IFC mod_2544 <- mkDebugOperation(mod_2544_inner, "mod_2544");
    Operation_IFC mod_2545_inner <- mkFlatten(2);
    Operation_IFC mod_2545 <- mkDebugOperation(mod_2545_inner, "mod_2545");
    Operation_IFC mod_2546_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2546 <- mkDebugOperation(mod_2546_inner, "mod_2546");
    Broadcast_IFC#(4) mod_2547_inner <- mkBroadcast(4);
    Operation_IFC mod_2547 <- mkDebugOperation(mod_2547_inner.op, "mod_2547");
    PMU_IFC mod_2548_bufferize <- mkPMU(2);
    Operation_IFC mod_2548_inner = mod_2548_bufferize.operation;
    Operation_IFC mod_2548 <- mkDebugOperation(mod_2548_inner, "mod_2548");
    Broadcast_IFC#(2) mod_2549_inner <- mkBroadcast(2);
    Operation_IFC mod_2549 <- mkDebugOperation(mod_2549_inner.op, "mod_2549");
    PMU_IFC mod_2550_bufferize <- mkPMU(1);
    Operation_IFC mod_2550_inner = mod_2550_bufferize.operation;
    Operation_IFC mod_2550 <- mkDebugOperation(mod_2550_inner, "mod_2550");
    Operation_IFC mod_2551_inner <- mkBinaryMap(1094, matmul_t_tile);
    Operation_IFC mod_2551 <- mkDebugOperation(mod_2551_inner, "mod_2551");
    Operation_IFC mod_2552_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2552 <- mkDebugOperation(mod_2552_inner, "mod_2552");
    Operation_IFC mod_2553_inner <- mkBinaryMap(1862, mul_tile);
    Operation_IFC mod_2553 <- mkDebugOperation(mod_2553_inner, "mod_2553");
    PMU_IFC mod_2554_bufferize <- mkPMU(1);
    Operation_IFC mod_2554_inner = mod_2554_bufferize.operation;
    Operation_IFC mod_2554 <- mkDebugOperation(mod_2554_inner, "mod_2554");
    Operation_IFC mod_2555_inner <- mkBinaryMap(2439, matmul_t_tile);
    Operation_IFC mod_2555 <- mkDebugOperation(mod_2555_inner, "mod_2555");
    Operation_IFC mod_2556_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2556 <- mkDebugOperation(mod_2556_inner, "mod_2556");
    Operation_IFC mod_2557_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2557 <- mkDebugOperation(mod_2557_inner, "mod_2557");
    Operation_IFC mod_2558_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2558 <- mkDebugOperation(mod_2558_inner, "mod_2558");
    Operation_IFC mod_2559_inner <- mkBinaryMap(2761, mul_tile);
    Operation_IFC mod_2559 <- mkDebugOperation(mod_2559_inner, "mod_2559");
    PMU_IFC mod_2560_bufferize <- mkPMU(1);
    Operation_IFC mod_2560_inner = mod_2560_bufferize.operation;
    Operation_IFC mod_2560 <- mkDebugOperation(mod_2560_inner, "mod_2560");
    PMU_IFC mod_2561_bufferize <- mkPMU(2);
    Operation_IFC mod_2561_inner = mod_2561_bufferize.operation;
    Operation_IFC mod_2561 <- mkDebugOperation(mod_2561_inner, "mod_2561");
    PMU_IFC mod_2562_bufferize <- mkPMU(2);
    Operation_IFC mod_2562_inner = mod_2562_bufferize.operation;
    Operation_IFC mod_2562 <- mkDebugOperation(mod_2562_inner, "mod_2562");
    Operation_IFC mod_2563_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2563 <- mkDebugOperation(mod_2563_inner, "mod_2563");
    Operation_IFC mod_2564_inner <- mkFlatten(1);
    Operation_IFC mod_2564 <- mkDebugOperation(mod_2564_inner, "mod_2564");
    Operation_IFC mod_2565_inner <- mkFlatten(0);
    Operation_IFC mod_2565 <- mkDebugOperation(mod_2565_inner, "mod_2565");
    Operation_IFC mod_2566_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2566 <- mkDebugOperation(mod_2566_inner, "mod_2566");
    Operation_IFC mod_2567_inner <- mkUnaryMap(1734, silu_tile);
    Operation_IFC mod_2567 <- mkDebugOperation(mod_2567_inner, "mod_2567");
    Operation_IFC mod_2568_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2568 <- mkDebugOperation(mod_2568_inner, "mod_2568");
    Operation_IFC mod_2569_inner <- mkBinaryMap(1606, matmul_t_tile);
    Operation_IFC mod_2569 <- mkDebugOperation(mod_2569_inner, "mod_2569");
    PMU_IFC mod_2570_bufferize <- mkPMU(2);
    Operation_IFC mod_2570_inner = mod_2570_bufferize.operation;
    Operation_IFC mod_2570 <- mkDebugOperation(mod_2570_inner, "mod_2570");
    Operation_IFC mod_2571_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2571 <- mkDebugOperation(mod_2571_inner, "mod_2571");
    Operation_IFC mod_2572_inner <- mkFlatten(1);
    Operation_IFC mod_2572 <- mkDebugOperation(mod_2572_inner, "mod_2572");
    Operation_IFC mod_2573_inner <- mkFlatten(0);
    Operation_IFC mod_2573 <- mkDebugOperation(mod_2573_inner, "mod_2573");
    PMU_IFC mod_2574_bufferize <- mkPMU(1);
    Operation_IFC mod_2574_inner = mod_2574_bufferize.operation;
    Operation_IFC mod_2574 <- mkDebugOperation(mod_2574_inner, "mod_2574");
    Operation_IFC mod_2575_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2575 <- mkDebugOperation(mod_2575_inner, "mod_2575");
    PMU_IFC mod_2576_bufferize <- mkPMU(2);
    Operation_IFC mod_2576_inner = mod_2576_bufferize.operation;
    Operation_IFC mod_2576 <- mkDebugOperation(mod_2576_inner, "mod_2576");
    Operation_IFC mod_2577_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2577 <- mkDebugOperation(mod_2577_inner, "mod_2577");
    Operation_IFC mod_2578_inner <- mkFlatten(1);
    Operation_IFC mod_2578 <- mkDebugOperation(mod_2578_inner, "mod_2578");
    Operation_IFC mod_2579_inner <- mkFlatten(0);
    Operation_IFC mod_2579 <- mkDebugOperation(mod_2579_inner, "mod_2579");
    Operation_IFC mod_2580_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2580 <- mkDebugOperation(mod_2580_inner, "mod_2580");
    Operation_IFC mod_2581_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2581 <- mkDebugOperation(mod_2581_inner, "mod_2581");
    PMU_IFC mod_2582_bufferize <- mkPMU(2);
    Operation_IFC mod_2582_inner = mod_2582_bufferize.operation;
    Operation_IFC mod_2582 <- mkDebugOperation(mod_2582_inner, "mod_2582");
    rule rule_3287;
        ChannelMessage t;
        t <- mod_2545.get(0);
        mod_2546.put(0, t);
    endrule
    rule rule_3288;
        ChannelMessage t;
        t <- mod_2549.get(1);
        mod_2550.put(0, t);
    endrule
    rule rule_3289;
        ChannelMessage t;
        t <- mod_2543.get(0);
        mod_2544.put(0, t);
    endrule
    rule rule_3290;
        ChannelMessage t;
        t <- mod_2560.get(1);
        mod_2558.put(1, t);
    endrule
    rule rule_3291;
        ChannelMessage t;
        t <- mod_2574.get(1);
        mod_2569.put(0, t);
    endrule
    rule rule_3292;
        ChannelMessage t;
        t <- mod_2567.get(0);
        mod_2553.put(1, t);
    endrule
    rule rule_3293;
        ChannelMessage t;
        t <- mod_2578.get(0);
        mod_2576.put(0, t);
    endrule
    rule rule_3294;
        ChannelMessage t;
        t <- mod_2582.get(0);
        mod_2582.put(1, t);
    endrule
    rule rule_3295;
        ChannelMessage t;
        t <- mod_2558.get(0);
        mod_2560.put(0, t);
    endrule
    rule rule_3296;
        ChannelMessage t;
        t <- mod_2547.get(3);
        mod_2548.put(0, t);
    endrule
    rule rule_3297;
        ChannelMessage t;
        t <- mod_2550.get(0);
        mod_2580.put(0, t);
    endrule
    rule rule_3298;
        ChannelMessage t;
        t <- mod_2581.get(0);
        mod_2548.put(1, t);
    endrule
    rule rule_3299;
        ChannelMessage t;
        t <- mod_2554.get(0);
        mod_2566.put(0, t);
    endrule
    rule rule_3300;
        ChannelMessage t;
        t <- mod_2548.get(1);
        mod_2549.put(0, t);
    endrule
    rule rule_3301;
        ChannelMessage t;
        t <- mod_2572.get(0);
        mod_2570.put(0, t);
    endrule
    rule rule_3302;
        ChannelMessage t;
        t <- mod_2548.get(0);
        mod_2581.put(0, t);
    endrule
    rule rule_3303;
        ChannelMessage t;
        t <- mod_2546.get(0);
        mod_2582.put(0, t);
    endrule
    rule rule_3304;
        ChannelMessage t;
        t <- mod_2557.get(1);
        mod_2558.put(0, t);
    endrule
    rule rule_3305;
        ChannelMessage t;
        t <- mod_2570.get(0);
        mod_2571.put(0, t);
    endrule
    rule rule_3306;
        ChannelMessage t;
        t <- mod_2566.get(0);
        mod_2554.put(1, t);
    endrule
    rule rule_3307;
        ChannelMessage t;
        t <- mod_2582.get(1);
        mod_2546.put(1, t);
    endrule
    rule rule_3308;
        ChannelMessage t;
        t <- mod_2577.get(0);
        mod_2576.put(1, t);
    endrule
    rule rule_3309;
        ChannelMessage t;
        t <- mod_2570.get(1);
        mod_2569.put(1, t);
    endrule
    rule rule_3310;
        ChannelMessage t;
        t <- mod_2555.get(0);
        mod_2556.put(0, t);
    endrule
    rule rule_3311;
        ChannelMessage t;
        t <- mod_2550.get(1);
        mod_2551.put(0, t);
    endrule
    rule rule_3312;
        ChannelMessage t;
        t <- mod_2579.get(0);
        mod_2578.put(0, t);
    endrule
    rule rule_3313;
        ChannelMessage t;
        t <- mod_2571.get(0);
        mod_2570.put(1, t);
    endrule
    rule rule_3314;
        ChannelMessage t;
        t <- mod_2568.get(0);
        mod_2567.put(0, t);
    endrule
    rule rule_3315;
        ChannelMessage t;
        t <- mod_2551.get(0);
        mod_2552.put(0, t);
    endrule
    rule rule_3316;
        ChannelMessage t;
        t <- mod_2564.get(0);
        mod_2562.put(0, t);
    endrule
    rule rule_3317;
        ChannelMessage t;
        t <- mod_2561.get(0);
        mod_2561.put(1, t);
    endrule
    rule rule_3318;
        ChannelMessage t;
        t <- mod_2563.get(0);
        mod_2562.put(1, t);
    endrule
    rule rule_3319;
        ChannelMessage t;
        t <- mod_2546.get(1);
        mod_2547.put(0, t);
    endrule
    rule rule_3320;
        ChannelMessage t;
        t <- mod_2573.get(0);
        mod_2572.put(0, t);
    endrule
    rule rule_3321;
        ChannelMessage t;
        t <- mod_2561.get(1);
        mod_2557.put(1, t);
    endrule
    rule rule_3322;
        ChannelMessage t;
        t <- mod_2576.get(1);
        mod_2551.put(1, t);
    endrule
    rule rule_3323;
        ChannelMessage t;
        t <- mod_2574.get(0);
        mod_2575.put(0, t);
    endrule
    rule rule_3324;
        ChannelMessage t;
        t <- mod_2560.get(0);
        mod_2560.put(1, t);
    endrule
    rule rule_3325;
        ChannelMessage t;
        t <- mod_2565.get(0);
        mod_2564.put(0, t);
    endrule
    rule rule_3326;
        ChannelMessage t;
        t <- mod_2556.get(0);
        mod_2557.put(0, t);
    endrule
    rule rule_3327;
        ChannelMessage t;
        t <- mod_2562.get(0);
        mod_2563.put(0, t);
    endrule
    rule rule_3328;
        ChannelMessage t;
        t <- mod_2553.get(0);
        mod_2554.put(0, t);
    endrule
    rule rule_3329;
        ChannelMessage t;
        t <- mod_2558.get(1);
        mod_2559.put(1, t);
    endrule
    rule rule_3330;
        ChannelMessage t;
        t <- mod_2569.get(0);
        mod_2568.put(0, t);
    endrule
    rule rule_3331;
        ChannelMessage t;
        t <- mod_2580.get(0);
        mod_2550.put(1, t);
    endrule
    rule rule_3332;
        ChannelMessage t;
        t <- mod_2575.get(0);
        mod_2574.put(1, t);
    endrule
    rule rule_3333;
        ChannelMessage t;
        t <- mod_2549.get(0);
        mod_2574.put(0, t);
    endrule
    rule rule_3334;
        ChannelMessage t;
        t <- mod_2552.get(0);
        mod_2553.put(0, t);
    endrule
    rule rule_3335;
        ChannelMessage t;
        t <- mod_2557.get(0);
        mod_2561.put(0, t);
    endrule
    rule rule_3336;
        ChannelMessage t;
        t <- mod_2544.get(0);
        mod_2545.put(0, t);
    endrule
    rule rule_3337;
        ChannelMessage t;
        t <- mod_2576.get(0);
        mod_2577.put(0, t);
    endrule
    rule rule_3338;
        ChannelMessage t;
        t <- mod_2554.get(1);
        mod_2555.put(0, t);
    endrule
    rule rule_3339;
        ChannelMessage t;
        t <- mod_2562.get(1);
        mod_2555.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2543.put(0, t);
        end
        if (i == 1) begin
            mod_2559.put(0, t);
        end
        if (i == 2) begin
            mod_2565.put(0, t);
        end
        if (i == 3) begin
            mod_2573.put(0, t);
        end
        if (i == 4) begin
            mod_2579.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_2547.get(0);
        end
        if (i == 3) begin
            t <- mod_2547.get(1);
        end
        if (i == 2) begin
            t <- mod_2547.get(2);
        end
        if (i == 1) begin
            t <- mod_2559.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6097 (Operation_IFC);
    Operation_IFC mod_2584_inner <- mkReshape(2, 64);
    Operation_IFC mod_2584 <- mkDebugOperation(mod_2584_inner, "mod_2584");
    Operation_IFC mod_2585_inner <- mkFlatten(1);
    Operation_IFC mod_2585 <- mkDebugOperation(mod_2585_inner, "mod_2585");
    Operation_IFC mod_2586_inner <- mkFlatten(2);
    Operation_IFC mod_2586 <- mkDebugOperation(mod_2586_inner, "mod_2586");
    Operation_IFC mod_2587_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2587 <- mkDebugOperation(mod_2587_inner, "mod_2587");
    Broadcast_IFC#(4) mod_2588_inner <- mkBroadcast(4);
    Operation_IFC mod_2588 <- mkDebugOperation(mod_2588_inner.op, "mod_2588");
    PMU_IFC mod_2589_bufferize <- mkPMU(2);
    Operation_IFC mod_2589_inner = mod_2589_bufferize.operation;
    Operation_IFC mod_2589 <- mkDebugOperation(mod_2589_inner, "mod_2589");
    Broadcast_IFC#(2) mod_2590_inner <- mkBroadcast(2);
    Operation_IFC mod_2590 <- mkDebugOperation(mod_2590_inner.op, "mod_2590");
    PMU_IFC mod_2591_bufferize <- mkPMU(1);
    Operation_IFC mod_2591_inner = mod_2591_bufferize.operation;
    Operation_IFC mod_2591 <- mkDebugOperation(mod_2591_inner, "mod_2591");
    Operation_IFC mod_2592_inner <- mkBinaryMap(1093, matmul_t_tile);
    Operation_IFC mod_2592 <- mkDebugOperation(mod_2592_inner, "mod_2592");
    Operation_IFC mod_2593_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2593 <- mkDebugOperation(mod_2593_inner, "mod_2593");
    Operation_IFC mod_2594_inner <- mkBinaryMap(1861, mul_tile);
    Operation_IFC mod_2594 <- mkDebugOperation(mod_2594_inner, "mod_2594");
    PMU_IFC mod_2595_bufferize <- mkPMU(1);
    Operation_IFC mod_2595_inner = mod_2595_bufferize.operation;
    Operation_IFC mod_2595 <- mkDebugOperation(mod_2595_inner, "mod_2595");
    Operation_IFC mod_2596_inner <- mkBinaryMap(2437, matmul_t_tile);
    Operation_IFC mod_2596 <- mkDebugOperation(mod_2596_inner, "mod_2596");
    Operation_IFC mod_2597_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2597 <- mkDebugOperation(mod_2597_inner, "mod_2597");
    Operation_IFC mod_2598_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2598 <- mkDebugOperation(mod_2598_inner, "mod_2598");
    Operation_IFC mod_2599_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2599 <- mkDebugOperation(mod_2599_inner, "mod_2599");
    Operation_IFC mod_2600_inner <- mkBinaryMap(2760, mul_tile);
    Operation_IFC mod_2600 <- mkDebugOperation(mod_2600_inner, "mod_2600");
    PMU_IFC mod_2601_bufferize <- mkPMU(1);
    Operation_IFC mod_2601_inner = mod_2601_bufferize.operation;
    Operation_IFC mod_2601 <- mkDebugOperation(mod_2601_inner, "mod_2601");
    PMU_IFC mod_2602_bufferize <- mkPMU(2);
    Operation_IFC mod_2602_inner = mod_2602_bufferize.operation;
    Operation_IFC mod_2602 <- mkDebugOperation(mod_2602_inner, "mod_2602");
    PMU_IFC mod_2603_bufferize <- mkPMU(2);
    Operation_IFC mod_2603_inner = mod_2603_bufferize.operation;
    Operation_IFC mod_2603 <- mkDebugOperation(mod_2603_inner, "mod_2603");
    Operation_IFC mod_2604_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2604 <- mkDebugOperation(mod_2604_inner, "mod_2604");
    Operation_IFC mod_2605_inner <- mkFlatten(1);
    Operation_IFC mod_2605 <- mkDebugOperation(mod_2605_inner, "mod_2605");
    Operation_IFC mod_2606_inner <- mkFlatten(0);
    Operation_IFC mod_2606 <- mkDebugOperation(mod_2606_inner, "mod_2606");
    Operation_IFC mod_2607_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2607 <- mkDebugOperation(mod_2607_inner, "mod_2607");
    Operation_IFC mod_2608_inner <- mkUnaryMap(1733, silu_tile);
    Operation_IFC mod_2608 <- mkDebugOperation(mod_2608_inner, "mod_2608");
    Operation_IFC mod_2609_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2609 <- mkDebugOperation(mod_2609_inner, "mod_2609");
    Operation_IFC mod_2610_inner <- mkBinaryMap(1605, matmul_t_tile);
    Operation_IFC mod_2610 <- mkDebugOperation(mod_2610_inner, "mod_2610");
    PMU_IFC mod_2611_bufferize <- mkPMU(2);
    Operation_IFC mod_2611_inner = mod_2611_bufferize.operation;
    Operation_IFC mod_2611 <- mkDebugOperation(mod_2611_inner, "mod_2611");
    Operation_IFC mod_2612_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2612 <- mkDebugOperation(mod_2612_inner, "mod_2612");
    Operation_IFC mod_2613_inner <- mkFlatten(1);
    Operation_IFC mod_2613 <- mkDebugOperation(mod_2613_inner, "mod_2613");
    Operation_IFC mod_2614_inner <- mkFlatten(0);
    Operation_IFC mod_2614 <- mkDebugOperation(mod_2614_inner, "mod_2614");
    PMU_IFC mod_2615_bufferize <- mkPMU(1);
    Operation_IFC mod_2615_inner = mod_2615_bufferize.operation;
    Operation_IFC mod_2615 <- mkDebugOperation(mod_2615_inner, "mod_2615");
    Operation_IFC mod_2616_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2616 <- mkDebugOperation(mod_2616_inner, "mod_2616");
    PMU_IFC mod_2617_bufferize <- mkPMU(2);
    Operation_IFC mod_2617_inner = mod_2617_bufferize.operation;
    Operation_IFC mod_2617 <- mkDebugOperation(mod_2617_inner, "mod_2617");
    Operation_IFC mod_2618_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2618 <- mkDebugOperation(mod_2618_inner, "mod_2618");
    Operation_IFC mod_2619_inner <- mkFlatten(1);
    Operation_IFC mod_2619 <- mkDebugOperation(mod_2619_inner, "mod_2619");
    Operation_IFC mod_2620_inner <- mkFlatten(0);
    Operation_IFC mod_2620 <- mkDebugOperation(mod_2620_inner, "mod_2620");
    Operation_IFC mod_2621_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2621 <- mkDebugOperation(mod_2621_inner, "mod_2621");
    Operation_IFC mod_2622_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2622 <- mkDebugOperation(mod_2622_inner, "mod_2622");
    PMU_IFC mod_2623_bufferize <- mkPMU(2);
    Operation_IFC mod_2623_inner = mod_2623_bufferize.operation;
    Operation_IFC mod_2623 <- mkDebugOperation(mod_2623_inner, "mod_2623");
    rule rule_3340;
        ChannelMessage t;
        t <- mod_2612.get(0);
        mod_2611.put(1, t);
    endrule
    rule rule_3341;
        ChannelMessage t;
        t <- mod_2616.get(0);
        mod_2615.put(1, t);
    endrule
    rule rule_3342;
        ChannelMessage t;
        t <- mod_2615.get(1);
        mod_2610.put(0, t);
    endrule
    rule rule_3343;
        ChannelMessage t;
        t <- mod_2584.get(0);
        mod_2585.put(0, t);
    endrule
    rule rule_3344;
        ChannelMessage t;
        t <- mod_2589.get(0);
        mod_2622.put(0, t);
    endrule
    rule rule_3345;
        ChannelMessage t;
        t <- mod_2589.get(1);
        mod_2590.put(0, t);
    endrule
    rule rule_3346;
        ChannelMessage t;
        t <- mod_2607.get(0);
        mod_2595.put(1, t);
    endrule
    rule rule_3347;
        ChannelMessage t;
        t <- mod_2590.get(1);
        mod_2591.put(0, t);
    endrule
    rule rule_3348;
        ChannelMessage t;
        t <- mod_2596.get(0);
        mod_2597.put(0, t);
    endrule
    rule rule_3349;
        ChannelMessage t;
        t <- mod_2598.get(0);
        mod_2602.put(0, t);
    endrule
    rule rule_3350;
        ChannelMessage t;
        t <- mod_2594.get(0);
        mod_2595.put(0, t);
    endrule
    rule rule_3351;
        ChannelMessage t;
        t <- mod_2587.get(1);
        mod_2588.put(0, t);
    endrule
    rule rule_3352;
        ChannelMessage t;
        t <- mod_2591.get(1);
        mod_2592.put(0, t);
    endrule
    rule rule_3353;
        ChannelMessage t;
        t <- mod_2618.get(0);
        mod_2617.put(1, t);
    endrule
    rule rule_3354;
        ChannelMessage t;
        t <- mod_2590.get(0);
        mod_2615.put(0, t);
    endrule
    rule rule_3355;
        ChannelMessage t;
        t <- mod_2620.get(0);
        mod_2619.put(0, t);
    endrule
    rule rule_3356;
        ChannelMessage t;
        t <- mod_2605.get(0);
        mod_2603.put(0, t);
    endrule
    rule rule_3357;
        ChannelMessage t;
        t <- mod_2588.get(3);
        mod_2589.put(0, t);
    endrule
    rule rule_3358;
        ChannelMessage t;
        t <- mod_2611.get(0);
        mod_2612.put(0, t);
    endrule
    rule rule_3359;
        ChannelMessage t;
        t <- mod_2585.get(0);
        mod_2586.put(0, t);
    endrule
    rule rule_3360;
        ChannelMessage t;
        t <- mod_2599.get(1);
        mod_2600.put(1, t);
    endrule
    rule rule_3361;
        ChannelMessage t;
        t <- mod_2621.get(0);
        mod_2591.put(1, t);
    endrule
    rule rule_3362;
        ChannelMessage t;
        t <- mod_2611.get(1);
        mod_2610.put(1, t);
    endrule
    rule rule_3363;
        ChannelMessage t;
        t <- mod_2613.get(0);
        mod_2611.put(0, t);
    endrule
    rule rule_3364;
        ChannelMessage t;
        t <- mod_2619.get(0);
        mod_2617.put(0, t);
    endrule
    rule rule_3365;
        ChannelMessage t;
        t <- mod_2610.get(0);
        mod_2609.put(0, t);
    endrule
    rule rule_3366;
        ChannelMessage t;
        t <- mod_2603.get(1);
        mod_2596.put(1, t);
    endrule
    rule rule_3367;
        ChannelMessage t;
        t <- mod_2604.get(0);
        mod_2603.put(1, t);
    endrule
    rule rule_3368;
        ChannelMessage t;
        t <- mod_2587.get(0);
        mod_2623.put(0, t);
    endrule
    rule rule_3369;
        ChannelMessage t;
        t <- mod_2595.get(1);
        mod_2596.put(0, t);
    endrule
    rule rule_3370;
        ChannelMessage t;
        t <- mod_2614.get(0);
        mod_2613.put(0, t);
    endrule
    rule rule_3371;
        ChannelMessage t;
        t <- mod_2622.get(0);
        mod_2589.put(1, t);
    endrule
    rule rule_3372;
        ChannelMessage t;
        t <- mod_2586.get(0);
        mod_2587.put(0, t);
    endrule
    rule rule_3373;
        ChannelMessage t;
        t <- mod_2608.get(0);
        mod_2594.put(1, t);
    endrule
    rule rule_3374;
        ChannelMessage t;
        t <- mod_2617.get(0);
        mod_2618.put(0, t);
    endrule
    rule rule_3375;
        ChannelMessage t;
        t <- mod_2592.get(0);
        mod_2593.put(0, t);
    endrule
    rule rule_3376;
        ChannelMessage t;
        t <- mod_2595.get(0);
        mod_2607.put(0, t);
    endrule
    rule rule_3377;
        ChannelMessage t;
        t <- mod_2606.get(0);
        mod_2605.put(0, t);
    endrule
    rule rule_3378;
        ChannelMessage t;
        t <- mod_2598.get(1);
        mod_2599.put(0, t);
    endrule
    rule rule_3379;
        ChannelMessage t;
        t <- mod_2609.get(0);
        mod_2608.put(0, t);
    endrule
    rule rule_3380;
        ChannelMessage t;
        t <- mod_2623.get(0);
        mod_2623.put(1, t);
    endrule
    rule rule_3381;
        ChannelMessage t;
        t <- mod_2593.get(0);
        mod_2594.put(0, t);
    endrule
    rule rule_3382;
        ChannelMessage t;
        t <- mod_2599.get(0);
        mod_2601.put(0, t);
    endrule
    rule rule_3383;
        ChannelMessage t;
        t <- mod_2603.get(0);
        mod_2604.put(0, t);
    endrule
    rule rule_3384;
        ChannelMessage t;
        t <- mod_2602.get(0);
        mod_2602.put(1, t);
    endrule
    rule rule_3385;
        ChannelMessage t;
        t <- mod_2597.get(0);
        mod_2598.put(0, t);
    endrule
    rule rule_3386;
        ChannelMessage t;
        t <- mod_2623.get(1);
        mod_2587.put(1, t);
    endrule
    rule rule_3387;
        ChannelMessage t;
        t <- mod_2615.get(0);
        mod_2616.put(0, t);
    endrule
    rule rule_3388;
        ChannelMessage t;
        t <- mod_2602.get(1);
        mod_2598.put(1, t);
    endrule
    rule rule_3389;
        ChannelMessage t;
        t <- mod_2601.get(0);
        mod_2601.put(1, t);
    endrule
    rule rule_3390;
        ChannelMessage t;
        t <- mod_2617.get(1);
        mod_2592.put(1, t);
    endrule
    rule rule_3391;
        ChannelMessage t;
        t <- mod_2601.get(1);
        mod_2599.put(1, t);
    endrule
    rule rule_3392;
        ChannelMessage t;
        t <- mod_2591.get(0);
        mod_2621.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2584.put(0, t);
        end
        if (i == 1) begin
            mod_2600.put(0, t);
        end
        if (i == 2) begin
            mod_2606.put(0, t);
        end
        if (i == 3) begin
            mod_2614.put(0, t);
        end
        if (i == 4) begin
            mod_2620.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_2588.get(0);
        end
        if (i == 2) begin
            t <- mod_2588.get(1);
        end
        if (i == 1) begin
            t <- mod_2588.get(2);
        end
        if (i == 3) begin
            t <- mod_2600.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6098 (Operation_IFC);
    Operation_IFC mod_2625_inner <- mkReshape(2, 64);
    Operation_IFC mod_2625 <- mkDebugOperation(mod_2625_inner, "mod_2625");
    Operation_IFC mod_2626_inner <- mkFlatten(1);
    Operation_IFC mod_2626 <- mkDebugOperation(mod_2626_inner, "mod_2626");
    Operation_IFC mod_2627_inner <- mkFlatten(2);
    Operation_IFC mod_2627 <- mkDebugOperation(mod_2627_inner, "mod_2627");
    Operation_IFC mod_2628_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2628 <- mkDebugOperation(mod_2628_inner, "mod_2628");
    Broadcast_IFC#(4) mod_2629_inner <- mkBroadcast(4);
    Operation_IFC mod_2629 <- mkDebugOperation(mod_2629_inner.op, "mod_2629");
    PMU_IFC mod_2630_bufferize <- mkPMU(2);
    Operation_IFC mod_2630_inner = mod_2630_bufferize.operation;
    Operation_IFC mod_2630 <- mkDebugOperation(mod_2630_inner, "mod_2630");
    Broadcast_IFC#(2) mod_2631_inner <- mkBroadcast(2);
    Operation_IFC mod_2631 <- mkDebugOperation(mod_2631_inner.op, "mod_2631");
    PMU_IFC mod_2632_bufferize <- mkPMU(1);
    Operation_IFC mod_2632_inner = mod_2632_bufferize.operation;
    Operation_IFC mod_2632 <- mkDebugOperation(mod_2632_inner, "mod_2632");
    Operation_IFC mod_2633_inner <- mkBinaryMap(1092, matmul_t_tile);
    Operation_IFC mod_2633 <- mkDebugOperation(mod_2633_inner, "mod_2633");
    Operation_IFC mod_2634_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2634 <- mkDebugOperation(mod_2634_inner, "mod_2634");
    Operation_IFC mod_2635_inner <- mkBinaryMap(1860, mul_tile);
    Operation_IFC mod_2635 <- mkDebugOperation(mod_2635_inner, "mod_2635");
    PMU_IFC mod_2636_bufferize <- mkPMU(1);
    Operation_IFC mod_2636_inner = mod_2636_bufferize.operation;
    Operation_IFC mod_2636 <- mkDebugOperation(mod_2636_inner, "mod_2636");
    Operation_IFC mod_2637_inner <- mkBinaryMap(2435, matmul_t_tile);
    Operation_IFC mod_2637 <- mkDebugOperation(mod_2637_inner, "mod_2637");
    Operation_IFC mod_2638_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2638 <- mkDebugOperation(mod_2638_inner, "mod_2638");
    Operation_IFC mod_2639_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2639 <- mkDebugOperation(mod_2639_inner, "mod_2639");
    Operation_IFC mod_2640_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2640 <- mkDebugOperation(mod_2640_inner, "mod_2640");
    Operation_IFC mod_2641_inner <- mkBinaryMap(2759, mul_tile);
    Operation_IFC mod_2641 <- mkDebugOperation(mod_2641_inner, "mod_2641");
    PMU_IFC mod_2642_bufferize <- mkPMU(1);
    Operation_IFC mod_2642_inner = mod_2642_bufferize.operation;
    Operation_IFC mod_2642 <- mkDebugOperation(mod_2642_inner, "mod_2642");
    PMU_IFC mod_2643_bufferize <- mkPMU(2);
    Operation_IFC mod_2643_inner = mod_2643_bufferize.operation;
    Operation_IFC mod_2643 <- mkDebugOperation(mod_2643_inner, "mod_2643");
    PMU_IFC mod_2644_bufferize <- mkPMU(2);
    Operation_IFC mod_2644_inner = mod_2644_bufferize.operation;
    Operation_IFC mod_2644 <- mkDebugOperation(mod_2644_inner, "mod_2644");
    Operation_IFC mod_2645_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2645 <- mkDebugOperation(mod_2645_inner, "mod_2645");
    Operation_IFC mod_2646_inner <- mkFlatten(1);
    Operation_IFC mod_2646 <- mkDebugOperation(mod_2646_inner, "mod_2646");
    Operation_IFC mod_2647_inner <- mkFlatten(0);
    Operation_IFC mod_2647 <- mkDebugOperation(mod_2647_inner, "mod_2647");
    Operation_IFC mod_2648_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2648 <- mkDebugOperation(mod_2648_inner, "mod_2648");
    Operation_IFC mod_2649_inner <- mkUnaryMap(1732, silu_tile);
    Operation_IFC mod_2649 <- mkDebugOperation(mod_2649_inner, "mod_2649");
    Operation_IFC mod_2650_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2650 <- mkDebugOperation(mod_2650_inner, "mod_2650");
    Operation_IFC mod_2651_inner <- mkBinaryMap(1604, matmul_t_tile);
    Operation_IFC mod_2651 <- mkDebugOperation(mod_2651_inner, "mod_2651");
    PMU_IFC mod_2652_bufferize <- mkPMU(2);
    Operation_IFC mod_2652_inner = mod_2652_bufferize.operation;
    Operation_IFC mod_2652 <- mkDebugOperation(mod_2652_inner, "mod_2652");
    Operation_IFC mod_2653_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2653 <- mkDebugOperation(mod_2653_inner, "mod_2653");
    Operation_IFC mod_2654_inner <- mkFlatten(1);
    Operation_IFC mod_2654 <- mkDebugOperation(mod_2654_inner, "mod_2654");
    Operation_IFC mod_2655_inner <- mkFlatten(0);
    Operation_IFC mod_2655 <- mkDebugOperation(mod_2655_inner, "mod_2655");
    PMU_IFC mod_2656_bufferize <- mkPMU(1);
    Operation_IFC mod_2656_inner = mod_2656_bufferize.operation;
    Operation_IFC mod_2656 <- mkDebugOperation(mod_2656_inner, "mod_2656");
    Operation_IFC mod_2657_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2657 <- mkDebugOperation(mod_2657_inner, "mod_2657");
    PMU_IFC mod_2658_bufferize <- mkPMU(2);
    Operation_IFC mod_2658_inner = mod_2658_bufferize.operation;
    Operation_IFC mod_2658 <- mkDebugOperation(mod_2658_inner, "mod_2658");
    Operation_IFC mod_2659_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2659 <- mkDebugOperation(mod_2659_inner, "mod_2659");
    Operation_IFC mod_2660_inner <- mkFlatten(1);
    Operation_IFC mod_2660 <- mkDebugOperation(mod_2660_inner, "mod_2660");
    Operation_IFC mod_2661_inner <- mkFlatten(0);
    Operation_IFC mod_2661 <- mkDebugOperation(mod_2661_inner, "mod_2661");
    Operation_IFC mod_2662_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2662 <- mkDebugOperation(mod_2662_inner, "mod_2662");
    Operation_IFC mod_2663_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2663 <- mkDebugOperation(mod_2663_inner, "mod_2663");
    PMU_IFC mod_2664_bufferize <- mkPMU(2);
    Operation_IFC mod_2664_inner = mod_2664_bufferize.operation;
    Operation_IFC mod_2664 <- mkDebugOperation(mod_2664_inner, "mod_2664");
    rule rule_3393;
        ChannelMessage t;
        t <- mod_2642.get(1);
        mod_2640.put(1, t);
    endrule
    rule rule_3394;
        ChannelMessage t;
        t <- mod_2629.get(3);
        mod_2630.put(0, t);
    endrule
    rule rule_3395;
        ChannelMessage t;
        t <- mod_2659.get(0);
        mod_2658.put(1, t);
    endrule
    rule rule_3396;
        ChannelMessage t;
        t <- mod_2633.get(0);
        mod_2634.put(0, t);
    endrule
    rule rule_3397;
        ChannelMessage t;
        t <- mod_2635.get(0);
        mod_2636.put(0, t);
    endrule
    rule rule_3398;
        ChannelMessage t;
        t <- mod_2656.get(1);
        mod_2651.put(0, t);
    endrule
    rule rule_3399;
        ChannelMessage t;
        t <- mod_2646.get(0);
        mod_2644.put(0, t);
    endrule
    rule rule_3400;
        ChannelMessage t;
        t <- mod_2652.get(0);
        mod_2653.put(0, t);
    endrule
    rule rule_3401;
        ChannelMessage t;
        t <- mod_2636.get(0);
        mod_2648.put(0, t);
    endrule
    rule rule_3402;
        ChannelMessage t;
        t <- mod_2644.get(0);
        mod_2645.put(0, t);
    endrule
    rule rule_3403;
        ChannelMessage t;
        t <- mod_2660.get(0);
        mod_2658.put(0, t);
    endrule
    rule rule_3404;
        ChannelMessage t;
        t <- mod_2636.get(1);
        mod_2637.put(0, t);
    endrule
    rule rule_3405;
        ChannelMessage t;
        t <- mod_2651.get(0);
        mod_2650.put(0, t);
    endrule
    rule rule_3406;
        ChannelMessage t;
        t <- mod_2627.get(0);
        mod_2628.put(0, t);
    endrule
    rule rule_3407;
        ChannelMessage t;
        t <- mod_2662.get(0);
        mod_2632.put(1, t);
    endrule
    rule rule_3408;
        ChannelMessage t;
        t <- mod_2643.get(0);
        mod_2643.put(1, t);
    endrule
    rule rule_3409;
        ChannelMessage t;
        t <- mod_2640.get(0);
        mod_2642.put(0, t);
    endrule
    rule rule_3410;
        ChannelMessage t;
        t <- mod_2661.get(0);
        mod_2660.put(0, t);
    endrule
    rule rule_3411;
        ChannelMessage t;
        t <- mod_2652.get(1);
        mod_2651.put(1, t);
    endrule
    rule rule_3412;
        ChannelMessage t;
        t <- mod_2648.get(0);
        mod_2636.put(1, t);
    endrule
    rule rule_3413;
        ChannelMessage t;
        t <- mod_2634.get(0);
        mod_2635.put(0, t);
    endrule
    rule rule_3414;
        ChannelMessage t;
        t <- mod_2625.get(0);
        mod_2626.put(0, t);
    endrule
    rule rule_3415;
        ChannelMessage t;
        t <- mod_2656.get(0);
        mod_2657.put(0, t);
    endrule
    rule rule_3416;
        ChannelMessage t;
        t <- mod_2626.get(0);
        mod_2627.put(0, t);
    endrule
    rule rule_3417;
        ChannelMessage t;
        t <- mod_2658.get(1);
        mod_2633.put(1, t);
    endrule
    rule rule_3418;
        ChannelMessage t;
        t <- mod_2631.get(0);
        mod_2656.put(0, t);
    endrule
    rule rule_3419;
        ChannelMessage t;
        t <- mod_2637.get(0);
        mod_2638.put(0, t);
    endrule
    rule rule_3420;
        ChannelMessage t;
        t <- mod_2640.get(1);
        mod_2641.put(1, t);
    endrule
    rule rule_3421;
        ChannelMessage t;
        t <- mod_2630.get(0);
        mod_2663.put(0, t);
    endrule
    rule rule_3422;
        ChannelMessage t;
        t <- mod_2631.get(1);
        mod_2632.put(0, t);
    endrule
    rule rule_3423;
        ChannelMessage t;
        t <- mod_2649.get(0);
        mod_2635.put(1, t);
    endrule
    rule rule_3424;
        ChannelMessage t;
        t <- mod_2632.get(0);
        mod_2662.put(0, t);
    endrule
    rule rule_3425;
        ChannelMessage t;
        t <- mod_2647.get(0);
        mod_2646.put(0, t);
    endrule
    rule rule_3426;
        ChannelMessage t;
        t <- mod_2664.get(1);
        mod_2628.put(1, t);
    endrule
    rule rule_3427;
        ChannelMessage t;
        t <- mod_2657.get(0);
        mod_2656.put(1, t);
    endrule
    rule rule_3428;
        ChannelMessage t;
        t <- mod_2654.get(0);
        mod_2652.put(0, t);
    endrule
    rule rule_3429;
        ChannelMessage t;
        t <- mod_2642.get(0);
        mod_2642.put(1, t);
    endrule
    rule rule_3430;
        ChannelMessage t;
        t <- mod_2650.get(0);
        mod_2649.put(0, t);
    endrule
    rule rule_3431;
        ChannelMessage t;
        t <- mod_2639.get(0);
        mod_2643.put(0, t);
    endrule
    rule rule_3432;
        ChannelMessage t;
        t <- mod_2639.get(1);
        mod_2640.put(0, t);
    endrule
    rule rule_3433;
        ChannelMessage t;
        t <- mod_2628.get(1);
        mod_2629.put(0, t);
    endrule
    rule rule_3434;
        ChannelMessage t;
        t <- mod_2653.get(0);
        mod_2652.put(1, t);
    endrule
    rule rule_3435;
        ChannelMessage t;
        t <- mod_2630.get(1);
        mod_2631.put(0, t);
    endrule
    rule rule_3436;
        ChannelMessage t;
        t <- mod_2628.get(0);
        mod_2664.put(0, t);
    endrule
    rule rule_3437;
        ChannelMessage t;
        t <- mod_2663.get(0);
        mod_2630.put(1, t);
    endrule
    rule rule_3438;
        ChannelMessage t;
        t <- mod_2638.get(0);
        mod_2639.put(0, t);
    endrule
    rule rule_3439;
        ChannelMessage t;
        t <- mod_2655.get(0);
        mod_2654.put(0, t);
    endrule
    rule rule_3440;
        ChannelMessage t;
        t <- mod_2658.get(0);
        mod_2659.put(0, t);
    endrule
    rule rule_3441;
        ChannelMessage t;
        t <- mod_2645.get(0);
        mod_2644.put(1, t);
    endrule
    rule rule_3442;
        ChannelMessage t;
        t <- mod_2644.get(1);
        mod_2637.put(1, t);
    endrule
    rule rule_3443;
        ChannelMessage t;
        t <- mod_2664.get(0);
        mod_2664.put(1, t);
    endrule
    rule rule_3444;
        ChannelMessage t;
        t <- mod_2632.get(1);
        mod_2633.put(0, t);
    endrule
    rule rule_3445;
        ChannelMessage t;
        t <- mod_2643.get(1);
        mod_2639.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2625.put(0, t);
        end
        if (i == 1) begin
            mod_2641.put(0, t);
        end
        if (i == 2) begin
            mod_2647.put(0, t);
        end
        if (i == 3) begin
            mod_2655.put(0, t);
        end
        if (i == 4) begin
            mod_2661.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 2) begin
            t <- mod_2629.get(0);
        end
        if (i == 0) begin
            t <- mod_2629.get(1);
        end
        if (i == 1) begin
            t <- mod_2629.get(2);
        end
        if (i == 3) begin
            t <- mod_2641.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6099 (Operation_IFC);
    Operation_IFC mod_2666_inner <- mkReshape(2, 64);
    Operation_IFC mod_2666 <- mkDebugOperation(mod_2666_inner, "mod_2666");
    Operation_IFC mod_2667_inner <- mkFlatten(1);
    Operation_IFC mod_2667 <- mkDebugOperation(mod_2667_inner, "mod_2667");
    Operation_IFC mod_2668_inner <- mkFlatten(2);
    Operation_IFC mod_2668 <- mkDebugOperation(mod_2668_inner, "mod_2668");
    Operation_IFC mod_2669_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2669 <- mkDebugOperation(mod_2669_inner, "mod_2669");
    Broadcast_IFC#(4) mod_2670_inner <- mkBroadcast(4);
    Operation_IFC mod_2670 <- mkDebugOperation(mod_2670_inner.op, "mod_2670");
    PMU_IFC mod_2671_bufferize <- mkPMU(2);
    Operation_IFC mod_2671_inner = mod_2671_bufferize.operation;
    Operation_IFC mod_2671 <- mkDebugOperation(mod_2671_inner, "mod_2671");
    Broadcast_IFC#(2) mod_2672_inner <- mkBroadcast(2);
    Operation_IFC mod_2672 <- mkDebugOperation(mod_2672_inner.op, "mod_2672");
    PMU_IFC mod_2673_bufferize <- mkPMU(1);
    Operation_IFC mod_2673_inner = mod_2673_bufferize.operation;
    Operation_IFC mod_2673 <- mkDebugOperation(mod_2673_inner, "mod_2673");
    Operation_IFC mod_2674_inner <- mkBinaryMap(1091, matmul_t_tile);
    Operation_IFC mod_2674 <- mkDebugOperation(mod_2674_inner, "mod_2674");
    Operation_IFC mod_2675_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2675 <- mkDebugOperation(mod_2675_inner, "mod_2675");
    Operation_IFC mod_2676_inner <- mkBinaryMap(1859, mul_tile);
    Operation_IFC mod_2676 <- mkDebugOperation(mod_2676_inner, "mod_2676");
    PMU_IFC mod_2677_bufferize <- mkPMU(1);
    Operation_IFC mod_2677_inner = mod_2677_bufferize.operation;
    Operation_IFC mod_2677 <- mkDebugOperation(mod_2677_inner, "mod_2677");
    Operation_IFC mod_2678_inner <- mkBinaryMap(2433, matmul_t_tile);
    Operation_IFC mod_2678 <- mkDebugOperation(mod_2678_inner, "mod_2678");
    Operation_IFC mod_2679_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2679 <- mkDebugOperation(mod_2679_inner, "mod_2679");
    Operation_IFC mod_2680_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2680 <- mkDebugOperation(mod_2680_inner, "mod_2680");
    Operation_IFC mod_2681_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2681 <- mkDebugOperation(mod_2681_inner, "mod_2681");
    Operation_IFC mod_2682_inner <- mkBinaryMap(2758, mul_tile);
    Operation_IFC mod_2682 <- mkDebugOperation(mod_2682_inner, "mod_2682");
    PMU_IFC mod_2683_bufferize <- mkPMU(1);
    Operation_IFC mod_2683_inner = mod_2683_bufferize.operation;
    Operation_IFC mod_2683 <- mkDebugOperation(mod_2683_inner, "mod_2683");
    PMU_IFC mod_2684_bufferize <- mkPMU(2);
    Operation_IFC mod_2684_inner = mod_2684_bufferize.operation;
    Operation_IFC mod_2684 <- mkDebugOperation(mod_2684_inner, "mod_2684");
    PMU_IFC mod_2685_bufferize <- mkPMU(2);
    Operation_IFC mod_2685_inner = mod_2685_bufferize.operation;
    Operation_IFC mod_2685 <- mkDebugOperation(mod_2685_inner, "mod_2685");
    Operation_IFC mod_2686_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2686 <- mkDebugOperation(mod_2686_inner, "mod_2686");
    Operation_IFC mod_2687_inner <- mkFlatten(1);
    Operation_IFC mod_2687 <- mkDebugOperation(mod_2687_inner, "mod_2687");
    Operation_IFC mod_2688_inner <- mkFlatten(0);
    Operation_IFC mod_2688 <- mkDebugOperation(mod_2688_inner, "mod_2688");
    Operation_IFC mod_2689_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2689 <- mkDebugOperation(mod_2689_inner, "mod_2689");
    Operation_IFC mod_2690_inner <- mkUnaryMap(1731, silu_tile);
    Operation_IFC mod_2690 <- mkDebugOperation(mod_2690_inner, "mod_2690");
    Operation_IFC mod_2691_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2691 <- mkDebugOperation(mod_2691_inner, "mod_2691");
    Operation_IFC mod_2692_inner <- mkBinaryMap(1603, matmul_t_tile);
    Operation_IFC mod_2692 <- mkDebugOperation(mod_2692_inner, "mod_2692");
    PMU_IFC mod_2693_bufferize <- mkPMU(2);
    Operation_IFC mod_2693_inner = mod_2693_bufferize.operation;
    Operation_IFC mod_2693 <- mkDebugOperation(mod_2693_inner, "mod_2693");
    Operation_IFC mod_2694_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2694 <- mkDebugOperation(mod_2694_inner, "mod_2694");
    Operation_IFC mod_2695_inner <- mkFlatten(1);
    Operation_IFC mod_2695 <- mkDebugOperation(mod_2695_inner, "mod_2695");
    Operation_IFC mod_2696_inner <- mkFlatten(0);
    Operation_IFC mod_2696 <- mkDebugOperation(mod_2696_inner, "mod_2696");
    PMU_IFC mod_2697_bufferize <- mkPMU(1);
    Operation_IFC mod_2697_inner = mod_2697_bufferize.operation;
    Operation_IFC mod_2697 <- mkDebugOperation(mod_2697_inner, "mod_2697");
    Operation_IFC mod_2698_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2698 <- mkDebugOperation(mod_2698_inner, "mod_2698");
    PMU_IFC mod_2699_bufferize <- mkPMU(2);
    Operation_IFC mod_2699_inner = mod_2699_bufferize.operation;
    Operation_IFC mod_2699 <- mkDebugOperation(mod_2699_inner, "mod_2699");
    Operation_IFC mod_2700_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2700 <- mkDebugOperation(mod_2700_inner, "mod_2700");
    Operation_IFC mod_2701_inner <- mkFlatten(1);
    Operation_IFC mod_2701 <- mkDebugOperation(mod_2701_inner, "mod_2701");
    Operation_IFC mod_2702_inner <- mkFlatten(0);
    Operation_IFC mod_2702 <- mkDebugOperation(mod_2702_inner, "mod_2702");
    Operation_IFC mod_2703_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2703 <- mkDebugOperation(mod_2703_inner, "mod_2703");
    Operation_IFC mod_2704_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2704 <- mkDebugOperation(mod_2704_inner, "mod_2704");
    PMU_IFC mod_2705_bufferize <- mkPMU(2);
    Operation_IFC mod_2705_inner = mod_2705_bufferize.operation;
    Operation_IFC mod_2705 <- mkDebugOperation(mod_2705_inner, "mod_2705");
    rule rule_3446;
        ChannelMessage t;
        t <- mod_2672.get(1);
        mod_2673.put(0, t);
    endrule
    rule rule_3447;
        ChannelMessage t;
        t <- mod_2681.get(1);
        mod_2682.put(1, t);
    endrule
    rule rule_3448;
        ChannelMessage t;
        t <- mod_2693.get(1);
        mod_2692.put(1, t);
    endrule
    rule rule_3449;
        ChannelMessage t;
        t <- mod_2683.get(1);
        mod_2681.put(1, t);
    endrule
    rule rule_3450;
        ChannelMessage t;
        t <- mod_2692.get(0);
        mod_2691.put(0, t);
    endrule
    rule rule_3451;
        ChannelMessage t;
        t <- mod_2677.get(0);
        mod_2689.put(0, t);
    endrule
    rule rule_3452;
        ChannelMessage t;
        t <- mod_2699.get(0);
        mod_2700.put(0, t);
    endrule
    rule rule_3453;
        ChannelMessage t;
        t <- mod_2675.get(0);
        mod_2676.put(0, t);
    endrule
    rule rule_3454;
        ChannelMessage t;
        t <- mod_2701.get(0);
        mod_2699.put(0, t);
    endrule
    rule rule_3455;
        ChannelMessage t;
        t <- mod_2705.get(1);
        mod_2669.put(1, t);
    endrule
    rule rule_3456;
        ChannelMessage t;
        t <- mod_2666.get(0);
        mod_2667.put(0, t);
    endrule
    rule rule_3457;
        ChannelMessage t;
        t <- mod_2693.get(0);
        mod_2694.put(0, t);
    endrule
    rule rule_3458;
        ChannelMessage t;
        t <- mod_2687.get(0);
        mod_2685.put(0, t);
    endrule
    rule rule_3459;
        ChannelMessage t;
        t <- mod_2686.get(0);
        mod_2685.put(1, t);
    endrule
    rule rule_3460;
        ChannelMessage t;
        t <- mod_2697.get(0);
        mod_2698.put(0, t);
    endrule
    rule rule_3461;
        ChannelMessage t;
        t <- mod_2699.get(1);
        mod_2674.put(1, t);
    endrule
    rule rule_3462;
        ChannelMessage t;
        t <- mod_2671.get(0);
        mod_2704.put(0, t);
    endrule
    rule rule_3463;
        ChannelMessage t;
        t <- mod_2674.get(0);
        mod_2675.put(0, t);
    endrule
    rule rule_3464;
        ChannelMessage t;
        t <- mod_2680.get(1);
        mod_2681.put(0, t);
    endrule
    rule rule_3465;
        ChannelMessage t;
        t <- mod_2694.get(0);
        mod_2693.put(1, t);
    endrule
    rule rule_3466;
        ChannelMessage t;
        t <- mod_2695.get(0);
        mod_2693.put(0, t);
    endrule
    rule rule_3467;
        ChannelMessage t;
        t <- mod_2704.get(0);
        mod_2671.put(1, t);
    endrule
    rule rule_3468;
        ChannelMessage t;
        t <- mod_2676.get(0);
        mod_2677.put(0, t);
    endrule
    rule rule_3469;
        ChannelMessage t;
        t <- mod_2685.get(1);
        mod_2678.put(1, t);
    endrule
    rule rule_3470;
        ChannelMessage t;
        t <- mod_2673.get(0);
        mod_2703.put(0, t);
    endrule
    rule rule_3471;
        ChannelMessage t;
        t <- mod_2700.get(0);
        mod_2699.put(1, t);
    endrule
    rule rule_3472;
        ChannelMessage t;
        t <- mod_2689.get(0);
        mod_2677.put(1, t);
    endrule
    rule rule_3473;
        ChannelMessage t;
        t <- mod_2684.get(0);
        mod_2684.put(1, t);
    endrule
    rule rule_3474;
        ChannelMessage t;
        t <- mod_2685.get(0);
        mod_2686.put(0, t);
    endrule
    rule rule_3475;
        ChannelMessage t;
        t <- mod_2678.get(0);
        mod_2679.put(0, t);
    endrule
    rule rule_3476;
        ChannelMessage t;
        t <- mod_2669.get(1);
        mod_2670.put(0, t);
    endrule
    rule rule_3477;
        ChannelMessage t;
        t <- mod_2698.get(0);
        mod_2697.put(1, t);
    endrule
    rule rule_3478;
        ChannelMessage t;
        t <- mod_2673.get(1);
        mod_2674.put(0, t);
    endrule
    rule rule_3479;
        ChannelMessage t;
        t <- mod_2688.get(0);
        mod_2687.put(0, t);
    endrule
    rule rule_3480;
        ChannelMessage t;
        t <- mod_2702.get(0);
        mod_2701.put(0, t);
    endrule
    rule rule_3481;
        ChannelMessage t;
        t <- mod_2668.get(0);
        mod_2669.put(0, t);
    endrule
    rule rule_3482;
        ChannelMessage t;
        t <- mod_2683.get(0);
        mod_2683.put(1, t);
    endrule
    rule rule_3483;
        ChannelMessage t;
        t <- mod_2669.get(0);
        mod_2705.put(0, t);
    endrule
    rule rule_3484;
        ChannelMessage t;
        t <- mod_2680.get(0);
        mod_2684.put(0, t);
    endrule
    rule rule_3485;
        ChannelMessage t;
        t <- mod_2696.get(0);
        mod_2695.put(0, t);
    endrule
    rule rule_3486;
        ChannelMessage t;
        t <- mod_2679.get(0);
        mod_2680.put(0, t);
    endrule
    rule rule_3487;
        ChannelMessage t;
        t <- mod_2703.get(0);
        mod_2673.put(1, t);
    endrule
    rule rule_3488;
        ChannelMessage t;
        t <- mod_2697.get(1);
        mod_2692.put(0, t);
    endrule
    rule rule_3489;
        ChannelMessage t;
        t <- mod_2705.get(0);
        mod_2705.put(1, t);
    endrule
    rule rule_3490;
        ChannelMessage t;
        t <- mod_2691.get(0);
        mod_2690.put(0, t);
    endrule
    rule rule_3491;
        ChannelMessage t;
        t <- mod_2677.get(1);
        mod_2678.put(0, t);
    endrule
    rule rule_3492;
        ChannelMessage t;
        t <- mod_2670.get(3);
        mod_2671.put(0, t);
    endrule
    rule rule_3493;
        ChannelMessage t;
        t <- mod_2681.get(0);
        mod_2683.put(0, t);
    endrule
    rule rule_3494;
        ChannelMessage t;
        t <- mod_2690.get(0);
        mod_2676.put(1, t);
    endrule
    rule rule_3495;
        ChannelMessage t;
        t <- mod_2667.get(0);
        mod_2668.put(0, t);
    endrule
    rule rule_3496;
        ChannelMessage t;
        t <- mod_2671.get(1);
        mod_2672.put(0, t);
    endrule
    rule rule_3497;
        ChannelMessage t;
        t <- mod_2672.get(0);
        mod_2697.put(0, t);
    endrule
    rule rule_3498;
        ChannelMessage t;
        t <- mod_2684.get(1);
        mod_2680.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2666.put(0, t);
        end
        if (i == 1) begin
            mod_2682.put(0, t);
        end
        if (i == 2) begin
            mod_2688.put(0, t);
        end
        if (i == 3) begin
            mod_2696.put(0, t);
        end
        if (i == 4) begin
            mod_2702.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_2670.get(0);
        end
        if (i == 2) begin
            t <- mod_2670.get(1);
        end
        if (i == 1) begin
            t <- mod_2670.get(2);
        end
        if (i == 0) begin
            t <- mod_2682.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6100 (Operation_IFC);
    Operation_IFC mod_2707_inner <- mkReshape(2, 64);
    Operation_IFC mod_2707 <- mkDebugOperation(mod_2707_inner, "mod_2707");
    Operation_IFC mod_2708_inner <- mkFlatten(1);
    Operation_IFC mod_2708 <- mkDebugOperation(mod_2708_inner, "mod_2708");
    Operation_IFC mod_2709_inner <- mkFlatten(2);
    Operation_IFC mod_2709 <- mkDebugOperation(mod_2709_inner, "mod_2709");
    Operation_IFC mod_2710_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2710 <- mkDebugOperation(mod_2710_inner, "mod_2710");
    Broadcast_IFC#(4) mod_2711_inner <- mkBroadcast(4);
    Operation_IFC mod_2711 <- mkDebugOperation(mod_2711_inner.op, "mod_2711");
    PMU_IFC mod_2712_bufferize <- mkPMU(2);
    Operation_IFC mod_2712_inner = mod_2712_bufferize.operation;
    Operation_IFC mod_2712 <- mkDebugOperation(mod_2712_inner, "mod_2712");
    Broadcast_IFC#(2) mod_2713_inner <- mkBroadcast(2);
    Operation_IFC mod_2713 <- mkDebugOperation(mod_2713_inner.op, "mod_2713");
    PMU_IFC mod_2714_bufferize <- mkPMU(1);
    Operation_IFC mod_2714_inner = mod_2714_bufferize.operation;
    Operation_IFC mod_2714 <- mkDebugOperation(mod_2714_inner, "mod_2714");
    Operation_IFC mod_2715_inner <- mkBinaryMap(1090, matmul_t_tile);
    Operation_IFC mod_2715 <- mkDebugOperation(mod_2715_inner, "mod_2715");
    Operation_IFC mod_2716_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2716 <- mkDebugOperation(mod_2716_inner, "mod_2716");
    Operation_IFC mod_2717_inner <- mkBinaryMap(1858, mul_tile);
    Operation_IFC mod_2717 <- mkDebugOperation(mod_2717_inner, "mod_2717");
    PMU_IFC mod_2718_bufferize <- mkPMU(1);
    Operation_IFC mod_2718_inner = mod_2718_bufferize.operation;
    Operation_IFC mod_2718 <- mkDebugOperation(mod_2718_inner, "mod_2718");
    Operation_IFC mod_2719_inner <- mkBinaryMap(2431, matmul_t_tile);
    Operation_IFC mod_2719 <- mkDebugOperation(mod_2719_inner, "mod_2719");
    Operation_IFC mod_2720_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2720 <- mkDebugOperation(mod_2720_inner, "mod_2720");
    Operation_IFC mod_2721_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2721 <- mkDebugOperation(mod_2721_inner, "mod_2721");
    Operation_IFC mod_2722_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2722 <- mkDebugOperation(mod_2722_inner, "mod_2722");
    Operation_IFC mod_2723_inner <- mkBinaryMap(2757, mul_tile);
    Operation_IFC mod_2723 <- mkDebugOperation(mod_2723_inner, "mod_2723");
    PMU_IFC mod_2724_bufferize <- mkPMU(1);
    Operation_IFC mod_2724_inner = mod_2724_bufferize.operation;
    Operation_IFC mod_2724 <- mkDebugOperation(mod_2724_inner, "mod_2724");
    PMU_IFC mod_2725_bufferize <- mkPMU(2);
    Operation_IFC mod_2725_inner = mod_2725_bufferize.operation;
    Operation_IFC mod_2725 <- mkDebugOperation(mod_2725_inner, "mod_2725");
    PMU_IFC mod_2726_bufferize <- mkPMU(2);
    Operation_IFC mod_2726_inner = mod_2726_bufferize.operation;
    Operation_IFC mod_2726 <- mkDebugOperation(mod_2726_inner, "mod_2726");
    Operation_IFC mod_2727_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2727 <- mkDebugOperation(mod_2727_inner, "mod_2727");
    Operation_IFC mod_2728_inner <- mkFlatten(1);
    Operation_IFC mod_2728 <- mkDebugOperation(mod_2728_inner, "mod_2728");
    Operation_IFC mod_2729_inner <- mkFlatten(0);
    Operation_IFC mod_2729 <- mkDebugOperation(mod_2729_inner, "mod_2729");
    Operation_IFC mod_2730_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2730 <- mkDebugOperation(mod_2730_inner, "mod_2730");
    Operation_IFC mod_2731_inner <- mkUnaryMap(1730, silu_tile);
    Operation_IFC mod_2731 <- mkDebugOperation(mod_2731_inner, "mod_2731");
    Operation_IFC mod_2732_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2732 <- mkDebugOperation(mod_2732_inner, "mod_2732");
    Operation_IFC mod_2733_inner <- mkBinaryMap(1602, matmul_t_tile);
    Operation_IFC mod_2733 <- mkDebugOperation(mod_2733_inner, "mod_2733");
    PMU_IFC mod_2734_bufferize <- mkPMU(2);
    Operation_IFC mod_2734_inner = mod_2734_bufferize.operation;
    Operation_IFC mod_2734 <- mkDebugOperation(mod_2734_inner, "mod_2734");
    Operation_IFC mod_2735_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2735 <- mkDebugOperation(mod_2735_inner, "mod_2735");
    Operation_IFC mod_2736_inner <- mkFlatten(1);
    Operation_IFC mod_2736 <- mkDebugOperation(mod_2736_inner, "mod_2736");
    Operation_IFC mod_2737_inner <- mkFlatten(0);
    Operation_IFC mod_2737 <- mkDebugOperation(mod_2737_inner, "mod_2737");
    PMU_IFC mod_2738_bufferize <- mkPMU(1);
    Operation_IFC mod_2738_inner = mod_2738_bufferize.operation;
    Operation_IFC mod_2738 <- mkDebugOperation(mod_2738_inner, "mod_2738");
    Operation_IFC mod_2739_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2739 <- mkDebugOperation(mod_2739_inner, "mod_2739");
    PMU_IFC mod_2740_bufferize <- mkPMU(2);
    Operation_IFC mod_2740_inner = mod_2740_bufferize.operation;
    Operation_IFC mod_2740 <- mkDebugOperation(mod_2740_inner, "mod_2740");
    Operation_IFC mod_2741_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2741 <- mkDebugOperation(mod_2741_inner, "mod_2741");
    Operation_IFC mod_2742_inner <- mkFlatten(1);
    Operation_IFC mod_2742 <- mkDebugOperation(mod_2742_inner, "mod_2742");
    Operation_IFC mod_2743_inner <- mkFlatten(0);
    Operation_IFC mod_2743 <- mkDebugOperation(mod_2743_inner, "mod_2743");
    Operation_IFC mod_2744_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2744 <- mkDebugOperation(mod_2744_inner, "mod_2744");
    Operation_IFC mod_2745_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2745 <- mkDebugOperation(mod_2745_inner, "mod_2745");
    PMU_IFC mod_2746_bufferize <- mkPMU(2);
    Operation_IFC mod_2746_inner = mod_2746_bufferize.operation;
    Operation_IFC mod_2746 <- mkDebugOperation(mod_2746_inner, "mod_2746");
    rule rule_3499;
        ChannelMessage t;
        t <- mod_2710.get(1);
        mod_2711.put(0, t);
    endrule
    rule rule_3500;
        ChannelMessage t;
        t <- mod_2722.get(1);
        mod_2723.put(1, t);
    endrule
    rule rule_3501;
        ChannelMessage t;
        t <- mod_2718.get(0);
        mod_2730.put(0, t);
    endrule
    rule rule_3502;
        ChannelMessage t;
        t <- mod_2738.get(1);
        mod_2733.put(0, t);
    endrule
    rule rule_3503;
        ChannelMessage t;
        t <- mod_2710.get(0);
        mod_2746.put(0, t);
    endrule
    rule rule_3504;
        ChannelMessage t;
        t <- mod_2716.get(0);
        mod_2717.put(0, t);
    endrule
    rule rule_3505;
        ChannelMessage t;
        t <- mod_2709.get(0);
        mod_2710.put(0, t);
    endrule
    rule rule_3506;
        ChannelMessage t;
        t <- mod_2724.get(0);
        mod_2724.put(1, t);
    endrule
    rule rule_3507;
        ChannelMessage t;
        t <- mod_2734.get(1);
        mod_2733.put(1, t);
    endrule
    rule rule_3508;
        ChannelMessage t;
        t <- mod_2736.get(0);
        mod_2734.put(0, t);
    endrule
    rule rule_3509;
        ChannelMessage t;
        t <- mod_2719.get(0);
        mod_2720.put(0, t);
    endrule
    rule rule_3510;
        ChannelMessage t;
        t <- mod_2714.get(0);
        mod_2744.put(0, t);
    endrule
    rule rule_3511;
        ChannelMessage t;
        t <- mod_2734.get(0);
        mod_2735.put(0, t);
    endrule
    rule rule_3512;
        ChannelMessage t;
        t <- mod_2713.get(0);
        mod_2738.put(0, t);
    endrule
    rule rule_3513;
        ChannelMessage t;
        t <- mod_2729.get(0);
        mod_2728.put(0, t);
    endrule
    rule rule_3514;
        ChannelMessage t;
        t <- mod_2738.get(0);
        mod_2739.put(0, t);
    endrule
    rule rule_3515;
        ChannelMessage t;
        t <- mod_2735.get(0);
        mod_2734.put(1, t);
    endrule
    rule rule_3516;
        ChannelMessage t;
        t <- mod_2711.get(3);
        mod_2712.put(0, t);
    endrule
    rule rule_3517;
        ChannelMessage t;
        t <- mod_2715.get(0);
        mod_2716.put(0, t);
    endrule
    rule rule_3518;
        ChannelMessage t;
        t <- mod_2726.get(1);
        mod_2719.put(1, t);
    endrule
    rule rule_3519;
        ChannelMessage t;
        t <- mod_2733.get(0);
        mod_2732.put(0, t);
    endrule
    rule rule_3520;
        ChannelMessage t;
        t <- mod_2713.get(1);
        mod_2714.put(0, t);
    endrule
    rule rule_3521;
        ChannelMessage t;
        t <- mod_2725.get(0);
        mod_2725.put(1, t);
    endrule
    rule rule_3522;
        ChannelMessage t;
        t <- mod_2708.get(0);
        mod_2709.put(0, t);
    endrule
    rule rule_3523;
        ChannelMessage t;
        t <- mod_2726.get(0);
        mod_2727.put(0, t);
    endrule
    rule rule_3524;
        ChannelMessage t;
        t <- mod_2721.get(0);
        mod_2725.put(0, t);
    endrule
    rule rule_3525;
        ChannelMessage t;
        t <- mod_2727.get(0);
        mod_2726.put(1, t);
    endrule
    rule rule_3526;
        ChannelMessage t;
        t <- mod_2740.get(0);
        mod_2741.put(0, t);
    endrule
    rule rule_3527;
        ChannelMessage t;
        t <- mod_2718.get(1);
        mod_2719.put(0, t);
    endrule
    rule rule_3528;
        ChannelMessage t;
        t <- mod_2746.get(0);
        mod_2746.put(1, t);
    endrule
    rule rule_3529;
        ChannelMessage t;
        t <- mod_2725.get(1);
        mod_2721.put(1, t);
    endrule
    rule rule_3530;
        ChannelMessage t;
        t <- mod_2740.get(1);
        mod_2715.put(1, t);
    endrule
    rule rule_3531;
        ChannelMessage t;
        t <- mod_2707.get(0);
        mod_2708.put(0, t);
    endrule
    rule rule_3532;
        ChannelMessage t;
        t <- mod_2724.get(1);
        mod_2722.put(1, t);
    endrule
    rule rule_3533;
        ChannelMessage t;
        t <- mod_2739.get(0);
        mod_2738.put(1, t);
    endrule
    rule rule_3534;
        ChannelMessage t;
        t <- mod_2742.get(0);
        mod_2740.put(0, t);
    endrule
    rule rule_3535;
        ChannelMessage t;
        t <- mod_2741.get(0);
        mod_2740.put(1, t);
    endrule
    rule rule_3536;
        ChannelMessage t;
        t <- mod_2714.get(1);
        mod_2715.put(0, t);
    endrule
    rule rule_3537;
        ChannelMessage t;
        t <- mod_2721.get(1);
        mod_2722.put(0, t);
    endrule
    rule rule_3538;
        ChannelMessage t;
        t <- mod_2744.get(0);
        mod_2714.put(1, t);
    endrule
    rule rule_3539;
        ChannelMessage t;
        t <- mod_2720.get(0);
        mod_2721.put(0, t);
    endrule
    rule rule_3540;
        ChannelMessage t;
        t <- mod_2712.get(0);
        mod_2745.put(0, t);
    endrule
    rule rule_3541;
        ChannelMessage t;
        t <- mod_2722.get(0);
        mod_2724.put(0, t);
    endrule
    rule rule_3542;
        ChannelMessage t;
        t <- mod_2728.get(0);
        mod_2726.put(0, t);
    endrule
    rule rule_3543;
        ChannelMessage t;
        t <- mod_2712.get(1);
        mod_2713.put(0, t);
    endrule
    rule rule_3544;
        ChannelMessage t;
        t <- mod_2717.get(0);
        mod_2718.put(0, t);
    endrule
    rule rule_3545;
        ChannelMessage t;
        t <- mod_2737.get(0);
        mod_2736.put(0, t);
    endrule
    rule rule_3546;
        ChannelMessage t;
        t <- mod_2731.get(0);
        mod_2717.put(1, t);
    endrule
    rule rule_3547;
        ChannelMessage t;
        t <- mod_2743.get(0);
        mod_2742.put(0, t);
    endrule
    rule rule_3548;
        ChannelMessage t;
        t <- mod_2745.get(0);
        mod_2712.put(1, t);
    endrule
    rule rule_3549;
        ChannelMessage t;
        t <- mod_2732.get(0);
        mod_2731.put(0, t);
    endrule
    rule rule_3550;
        ChannelMessage t;
        t <- mod_2730.get(0);
        mod_2718.put(1, t);
    endrule
    rule rule_3551;
        ChannelMessage t;
        t <- mod_2746.get(1);
        mod_2710.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2707.put(0, t);
        end
        if (i == 1) begin
            mod_2723.put(0, t);
        end
        if (i == 2) begin
            mod_2729.put(0, t);
        end
        if (i == 3) begin
            mod_2737.put(0, t);
        end
        if (i == 4) begin
            mod_2743.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_2711.get(0);
        end
        if (i == 3) begin
            t <- mod_2711.get(1);
        end
        if (i == 2) begin
            t <- mod_2711.get(2);
        end
        if (i == 1) begin
            t <- mod_2723.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6101 (Operation_IFC);
    Operation_IFC mod_2748_inner <- mkReshape(2, 64);
    Operation_IFC mod_2748 <- mkDebugOperation(mod_2748_inner, "mod_2748");
    Operation_IFC mod_2749_inner <- mkFlatten(1);
    Operation_IFC mod_2749 <- mkDebugOperation(mod_2749_inner, "mod_2749");
    Operation_IFC mod_2750_inner <- mkFlatten(2);
    Operation_IFC mod_2750 <- mkDebugOperation(mod_2750_inner, "mod_2750");
    Operation_IFC mod_2751_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2751 <- mkDebugOperation(mod_2751_inner, "mod_2751");
    Broadcast_IFC#(4) mod_2752_inner <- mkBroadcast(4);
    Operation_IFC mod_2752 <- mkDebugOperation(mod_2752_inner.op, "mod_2752");
    PMU_IFC mod_2753_bufferize <- mkPMU(2);
    Operation_IFC mod_2753_inner = mod_2753_bufferize.operation;
    Operation_IFC mod_2753 <- mkDebugOperation(mod_2753_inner, "mod_2753");
    Broadcast_IFC#(2) mod_2754_inner <- mkBroadcast(2);
    Operation_IFC mod_2754 <- mkDebugOperation(mod_2754_inner.op, "mod_2754");
    PMU_IFC mod_2755_bufferize <- mkPMU(1);
    Operation_IFC mod_2755_inner = mod_2755_bufferize.operation;
    Operation_IFC mod_2755 <- mkDebugOperation(mod_2755_inner, "mod_2755");
    Operation_IFC mod_2756_inner <- mkBinaryMap(1089, matmul_t_tile);
    Operation_IFC mod_2756 <- mkDebugOperation(mod_2756_inner, "mod_2756");
    Operation_IFC mod_2757_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2757 <- mkDebugOperation(mod_2757_inner, "mod_2757");
    Operation_IFC mod_2758_inner <- mkBinaryMap(1857, mul_tile);
    Operation_IFC mod_2758 <- mkDebugOperation(mod_2758_inner, "mod_2758");
    PMU_IFC mod_2759_bufferize <- mkPMU(1);
    Operation_IFC mod_2759_inner = mod_2759_bufferize.operation;
    Operation_IFC mod_2759 <- mkDebugOperation(mod_2759_inner, "mod_2759");
    Operation_IFC mod_2760_inner <- mkBinaryMap(2429, matmul_t_tile);
    Operation_IFC mod_2760 <- mkDebugOperation(mod_2760_inner, "mod_2760");
    Operation_IFC mod_2761_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2761 <- mkDebugOperation(mod_2761_inner, "mod_2761");
    Operation_IFC mod_2762_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2762 <- mkDebugOperation(mod_2762_inner, "mod_2762");
    Operation_IFC mod_2763_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2763 <- mkDebugOperation(mod_2763_inner, "mod_2763");
    Operation_IFC mod_2764_inner <- mkBinaryMap(2756, mul_tile);
    Operation_IFC mod_2764 <- mkDebugOperation(mod_2764_inner, "mod_2764");
    PMU_IFC mod_2765_bufferize <- mkPMU(1);
    Operation_IFC mod_2765_inner = mod_2765_bufferize.operation;
    Operation_IFC mod_2765 <- mkDebugOperation(mod_2765_inner, "mod_2765");
    PMU_IFC mod_2766_bufferize <- mkPMU(2);
    Operation_IFC mod_2766_inner = mod_2766_bufferize.operation;
    Operation_IFC mod_2766 <- mkDebugOperation(mod_2766_inner, "mod_2766");
    PMU_IFC mod_2767_bufferize <- mkPMU(2);
    Operation_IFC mod_2767_inner = mod_2767_bufferize.operation;
    Operation_IFC mod_2767 <- mkDebugOperation(mod_2767_inner, "mod_2767");
    Operation_IFC mod_2768_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2768 <- mkDebugOperation(mod_2768_inner, "mod_2768");
    Operation_IFC mod_2769_inner <- mkFlatten(1);
    Operation_IFC mod_2769 <- mkDebugOperation(mod_2769_inner, "mod_2769");
    Operation_IFC mod_2770_inner <- mkFlatten(0);
    Operation_IFC mod_2770 <- mkDebugOperation(mod_2770_inner, "mod_2770");
    Operation_IFC mod_2771_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2771 <- mkDebugOperation(mod_2771_inner, "mod_2771");
    Operation_IFC mod_2772_inner <- mkUnaryMap(1729, silu_tile);
    Operation_IFC mod_2772 <- mkDebugOperation(mod_2772_inner, "mod_2772");
    Operation_IFC mod_2773_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2773 <- mkDebugOperation(mod_2773_inner, "mod_2773");
    Operation_IFC mod_2774_inner <- mkBinaryMap(1601, matmul_t_tile);
    Operation_IFC mod_2774 <- mkDebugOperation(mod_2774_inner, "mod_2774");
    PMU_IFC mod_2775_bufferize <- mkPMU(2);
    Operation_IFC mod_2775_inner = mod_2775_bufferize.operation;
    Operation_IFC mod_2775 <- mkDebugOperation(mod_2775_inner, "mod_2775");
    Operation_IFC mod_2776_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2776 <- mkDebugOperation(mod_2776_inner, "mod_2776");
    Operation_IFC mod_2777_inner <- mkFlatten(1);
    Operation_IFC mod_2777 <- mkDebugOperation(mod_2777_inner, "mod_2777");
    Operation_IFC mod_2778_inner <- mkFlatten(0);
    Operation_IFC mod_2778 <- mkDebugOperation(mod_2778_inner, "mod_2778");
    PMU_IFC mod_2779_bufferize <- mkPMU(1);
    Operation_IFC mod_2779_inner = mod_2779_bufferize.operation;
    Operation_IFC mod_2779 <- mkDebugOperation(mod_2779_inner, "mod_2779");
    Operation_IFC mod_2780_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2780 <- mkDebugOperation(mod_2780_inner, "mod_2780");
    PMU_IFC mod_2781_bufferize <- mkPMU(2);
    Operation_IFC mod_2781_inner = mod_2781_bufferize.operation;
    Operation_IFC mod_2781 <- mkDebugOperation(mod_2781_inner, "mod_2781");
    Operation_IFC mod_2782_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2782 <- mkDebugOperation(mod_2782_inner, "mod_2782");
    Operation_IFC mod_2783_inner <- mkFlatten(1);
    Operation_IFC mod_2783 <- mkDebugOperation(mod_2783_inner, "mod_2783");
    Operation_IFC mod_2784_inner <- mkFlatten(0);
    Operation_IFC mod_2784 <- mkDebugOperation(mod_2784_inner, "mod_2784");
    Operation_IFC mod_2785_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2785 <- mkDebugOperation(mod_2785_inner, "mod_2785");
    Operation_IFC mod_2786_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2786 <- mkDebugOperation(mod_2786_inner, "mod_2786");
    PMU_IFC mod_2787_bufferize <- mkPMU(2);
    Operation_IFC mod_2787_inner = mod_2787_bufferize.operation;
    Operation_IFC mod_2787 <- mkDebugOperation(mod_2787_inner, "mod_2787");
    rule rule_3552;
        ChannelMessage t;
        t <- mod_2752.get(3);
        mod_2753.put(0, t);
    endrule
    rule rule_3553;
        ChannelMessage t;
        t <- mod_2769.get(0);
        mod_2767.put(0, t);
    endrule
    rule rule_3554;
        ChannelMessage t;
        t <- mod_2770.get(0);
        mod_2769.put(0, t);
    endrule
    rule rule_3555;
        ChannelMessage t;
        t <- mod_2754.get(0);
        mod_2779.put(0, t);
    endrule
    rule rule_3556;
        ChannelMessage t;
        t <- mod_2774.get(0);
        mod_2773.put(0, t);
    endrule
    rule rule_3557;
        ChannelMessage t;
        t <- mod_2780.get(0);
        mod_2779.put(1, t);
    endrule
    rule rule_3558;
        ChannelMessage t;
        t <- mod_2750.get(0);
        mod_2751.put(0, t);
    endrule
    rule rule_3559;
        ChannelMessage t;
        t <- mod_2751.get(0);
        mod_2787.put(0, t);
    endrule
    rule rule_3560;
        ChannelMessage t;
        t <- mod_2761.get(0);
        mod_2762.put(0, t);
    endrule
    rule rule_3561;
        ChannelMessage t;
        t <- mod_2787.get(1);
        mod_2751.put(1, t);
    endrule
    rule rule_3562;
        ChannelMessage t;
        t <- mod_2759.get(0);
        mod_2771.put(0, t);
    endrule
    rule rule_3563;
        ChannelMessage t;
        t <- mod_2779.get(0);
        mod_2780.put(0, t);
    endrule
    rule rule_3564;
        ChannelMessage t;
        t <- mod_2748.get(0);
        mod_2749.put(0, t);
    endrule
    rule rule_3565;
        ChannelMessage t;
        t <- mod_2766.get(1);
        mod_2762.put(1, t);
    endrule
    rule rule_3566;
        ChannelMessage t;
        t <- mod_2786.get(0);
        mod_2753.put(1, t);
    endrule
    rule rule_3567;
        ChannelMessage t;
        t <- mod_2775.get(1);
        mod_2774.put(1, t);
    endrule
    rule rule_3568;
        ChannelMessage t;
        t <- mod_2777.get(0);
        mod_2775.put(0, t);
    endrule
    rule rule_3569;
        ChannelMessage t;
        t <- mod_2763.get(1);
        mod_2764.put(1, t);
    endrule
    rule rule_3570;
        ChannelMessage t;
        t <- mod_2787.get(0);
        mod_2787.put(1, t);
    endrule
    rule rule_3571;
        ChannelMessage t;
        t <- mod_2758.get(0);
        mod_2759.put(0, t);
    endrule
    rule rule_3572;
        ChannelMessage t;
        t <- mod_2751.get(1);
        mod_2752.put(0, t);
    endrule
    rule rule_3573;
        ChannelMessage t;
        t <- mod_2767.get(1);
        mod_2760.put(1, t);
    endrule
    rule rule_3574;
        ChannelMessage t;
        t <- mod_2785.get(0);
        mod_2755.put(1, t);
    endrule
    rule rule_3575;
        ChannelMessage t;
        t <- mod_2754.get(1);
        mod_2755.put(0, t);
    endrule
    rule rule_3576;
        ChannelMessage t;
        t <- mod_2757.get(0);
        mod_2758.put(0, t);
    endrule
    rule rule_3577;
        ChannelMessage t;
        t <- mod_2784.get(0);
        mod_2783.put(0, t);
    endrule
    rule rule_3578;
        ChannelMessage t;
        t <- mod_2762.get(0);
        mod_2766.put(0, t);
    endrule
    rule rule_3579;
        ChannelMessage t;
        t <- mod_2779.get(1);
        mod_2774.put(0, t);
    endrule
    rule rule_3580;
        ChannelMessage t;
        t <- mod_2781.get(1);
        mod_2756.put(1, t);
    endrule
    rule rule_3581;
        ChannelMessage t;
        t <- mod_2765.get(0);
        mod_2765.put(1, t);
    endrule
    rule rule_3582;
        ChannelMessage t;
        t <- mod_2767.get(0);
        mod_2768.put(0, t);
    endrule
    rule rule_3583;
        ChannelMessage t;
        t <- mod_2772.get(0);
        mod_2758.put(1, t);
    endrule
    rule rule_3584;
        ChannelMessage t;
        t <- mod_2778.get(0);
        mod_2777.put(0, t);
    endrule
    rule rule_3585;
        ChannelMessage t;
        t <- mod_2749.get(0);
        mod_2750.put(0, t);
    endrule
    rule rule_3586;
        ChannelMessage t;
        t <- mod_2753.get(0);
        mod_2786.put(0, t);
    endrule
    rule rule_3587;
        ChannelMessage t;
        t <- mod_2762.get(1);
        mod_2763.put(0, t);
    endrule
    rule rule_3588;
        ChannelMessage t;
        t <- mod_2775.get(0);
        mod_2776.put(0, t);
    endrule
    rule rule_3589;
        ChannelMessage t;
        t <- mod_2783.get(0);
        mod_2781.put(0, t);
    endrule
    rule rule_3590;
        ChannelMessage t;
        t <- mod_2756.get(0);
        mod_2757.put(0, t);
    endrule
    rule rule_3591;
        ChannelMessage t;
        t <- mod_2766.get(0);
        mod_2766.put(1, t);
    endrule
    rule rule_3592;
        ChannelMessage t;
        t <- mod_2755.get(1);
        mod_2756.put(0, t);
    endrule
    rule rule_3593;
        ChannelMessage t;
        t <- mod_2765.get(1);
        mod_2763.put(1, t);
    endrule
    rule rule_3594;
        ChannelMessage t;
        t <- mod_2768.get(0);
        mod_2767.put(1, t);
    endrule
    rule rule_3595;
        ChannelMessage t;
        t <- mod_2773.get(0);
        mod_2772.put(0, t);
    endrule
    rule rule_3596;
        ChannelMessage t;
        t <- mod_2763.get(0);
        mod_2765.put(0, t);
    endrule
    rule rule_3597;
        ChannelMessage t;
        t <- mod_2781.get(0);
        mod_2782.put(0, t);
    endrule
    rule rule_3598;
        ChannelMessage t;
        t <- mod_2759.get(1);
        mod_2760.put(0, t);
    endrule
    rule rule_3599;
        ChannelMessage t;
        t <- mod_2753.get(1);
        mod_2754.put(0, t);
    endrule
    rule rule_3600;
        ChannelMessage t;
        t <- mod_2755.get(0);
        mod_2785.put(0, t);
    endrule
    rule rule_3601;
        ChannelMessage t;
        t <- mod_2771.get(0);
        mod_2759.put(1, t);
    endrule
    rule rule_3602;
        ChannelMessage t;
        t <- mod_2776.get(0);
        mod_2775.put(1, t);
    endrule
    rule rule_3603;
        ChannelMessage t;
        t <- mod_2782.get(0);
        mod_2781.put(1, t);
    endrule
    rule rule_3604;
        ChannelMessage t;
        t <- mod_2760.get(0);
        mod_2761.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2748.put(0, t);
        end
        if (i == 1) begin
            mod_2764.put(0, t);
        end
        if (i == 2) begin
            mod_2770.put(0, t);
        end
        if (i == 3) begin
            mod_2778.put(0, t);
        end
        if (i == 4) begin
            mod_2784.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_2752.get(0);
        end
        if (i == 3) begin
            t <- mod_2752.get(1);
        end
        if (i == 0) begin
            t <- mod_2752.get(2);
        end
        if (i == 2) begin
            t <- mod_2764.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6102 (Operation_IFC);
    Operation_IFC mod_2789_inner <- mkReshape(2, 64);
    Operation_IFC mod_2789 <- mkDebugOperation(mod_2789_inner, "mod_2789");
    Operation_IFC mod_2790_inner <- mkFlatten(1);
    Operation_IFC mod_2790 <- mkDebugOperation(mod_2790_inner, "mod_2790");
    Operation_IFC mod_2791_inner <- mkFlatten(2);
    Operation_IFC mod_2791 <- mkDebugOperation(mod_2791_inner, "mod_2791");
    Operation_IFC mod_2792_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2792 <- mkDebugOperation(mod_2792_inner, "mod_2792");
    Broadcast_IFC#(4) mod_2793_inner <- mkBroadcast(4);
    Operation_IFC mod_2793 <- mkDebugOperation(mod_2793_inner.op, "mod_2793");
    PMU_IFC mod_2794_bufferize <- mkPMU(2);
    Operation_IFC mod_2794_inner = mod_2794_bufferize.operation;
    Operation_IFC mod_2794 <- mkDebugOperation(mod_2794_inner, "mod_2794");
    Broadcast_IFC#(2) mod_2795_inner <- mkBroadcast(2);
    Operation_IFC mod_2795 <- mkDebugOperation(mod_2795_inner.op, "mod_2795");
    PMU_IFC mod_2796_bufferize <- mkPMU(1);
    Operation_IFC mod_2796_inner = mod_2796_bufferize.operation;
    Operation_IFC mod_2796 <- mkDebugOperation(mod_2796_inner, "mod_2796");
    Operation_IFC mod_2797_inner <- mkBinaryMap(1088, matmul_t_tile);
    Operation_IFC mod_2797 <- mkDebugOperation(mod_2797_inner, "mod_2797");
    Operation_IFC mod_2798_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2798 <- mkDebugOperation(mod_2798_inner, "mod_2798");
    Operation_IFC mod_2799_inner <- mkBinaryMap(1856, mul_tile);
    Operation_IFC mod_2799 <- mkDebugOperation(mod_2799_inner, "mod_2799");
    PMU_IFC mod_2800_bufferize <- mkPMU(1);
    Operation_IFC mod_2800_inner = mod_2800_bufferize.operation;
    Operation_IFC mod_2800 <- mkDebugOperation(mod_2800_inner, "mod_2800");
    Operation_IFC mod_2801_inner <- mkBinaryMap(2427, matmul_t_tile);
    Operation_IFC mod_2801 <- mkDebugOperation(mod_2801_inner, "mod_2801");
    Operation_IFC mod_2802_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2802 <- mkDebugOperation(mod_2802_inner, "mod_2802");
    Operation_IFC mod_2803_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2803 <- mkDebugOperation(mod_2803_inner, "mod_2803");
    Operation_IFC mod_2804_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2804 <- mkDebugOperation(mod_2804_inner, "mod_2804");
    Operation_IFC mod_2805_inner <- mkBinaryMap(2755, mul_tile);
    Operation_IFC mod_2805 <- mkDebugOperation(mod_2805_inner, "mod_2805");
    PMU_IFC mod_2806_bufferize <- mkPMU(1);
    Operation_IFC mod_2806_inner = mod_2806_bufferize.operation;
    Operation_IFC mod_2806 <- mkDebugOperation(mod_2806_inner, "mod_2806");
    PMU_IFC mod_2807_bufferize <- mkPMU(2);
    Operation_IFC mod_2807_inner = mod_2807_bufferize.operation;
    Operation_IFC mod_2807 <- mkDebugOperation(mod_2807_inner, "mod_2807");
    PMU_IFC mod_2808_bufferize <- mkPMU(2);
    Operation_IFC mod_2808_inner = mod_2808_bufferize.operation;
    Operation_IFC mod_2808 <- mkDebugOperation(mod_2808_inner, "mod_2808");
    Operation_IFC mod_2809_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2809 <- mkDebugOperation(mod_2809_inner, "mod_2809");
    Operation_IFC mod_2810_inner <- mkFlatten(1);
    Operation_IFC mod_2810 <- mkDebugOperation(mod_2810_inner, "mod_2810");
    Operation_IFC mod_2811_inner <- mkFlatten(0);
    Operation_IFC mod_2811 <- mkDebugOperation(mod_2811_inner, "mod_2811");
    Operation_IFC mod_2812_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2812 <- mkDebugOperation(mod_2812_inner, "mod_2812");
    Operation_IFC mod_2813_inner <- mkUnaryMap(1728, silu_tile);
    Operation_IFC mod_2813 <- mkDebugOperation(mod_2813_inner, "mod_2813");
    Operation_IFC mod_2814_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2814 <- mkDebugOperation(mod_2814_inner, "mod_2814");
    Operation_IFC mod_2815_inner <- mkBinaryMap(1600, matmul_t_tile);
    Operation_IFC mod_2815 <- mkDebugOperation(mod_2815_inner, "mod_2815");
    PMU_IFC mod_2816_bufferize <- mkPMU(2);
    Operation_IFC mod_2816_inner = mod_2816_bufferize.operation;
    Operation_IFC mod_2816 <- mkDebugOperation(mod_2816_inner, "mod_2816");
    Operation_IFC mod_2817_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2817 <- mkDebugOperation(mod_2817_inner, "mod_2817");
    Operation_IFC mod_2818_inner <- mkFlatten(1);
    Operation_IFC mod_2818 <- mkDebugOperation(mod_2818_inner, "mod_2818");
    Operation_IFC mod_2819_inner <- mkFlatten(0);
    Operation_IFC mod_2819 <- mkDebugOperation(mod_2819_inner, "mod_2819");
    PMU_IFC mod_2820_bufferize <- mkPMU(1);
    Operation_IFC mod_2820_inner = mod_2820_bufferize.operation;
    Operation_IFC mod_2820 <- mkDebugOperation(mod_2820_inner, "mod_2820");
    Operation_IFC mod_2821_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2821 <- mkDebugOperation(mod_2821_inner, "mod_2821");
    PMU_IFC mod_2822_bufferize <- mkPMU(2);
    Operation_IFC mod_2822_inner = mod_2822_bufferize.operation;
    Operation_IFC mod_2822 <- mkDebugOperation(mod_2822_inner, "mod_2822");
    Operation_IFC mod_2823_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2823 <- mkDebugOperation(mod_2823_inner, "mod_2823");
    Operation_IFC mod_2824_inner <- mkFlatten(1);
    Operation_IFC mod_2824 <- mkDebugOperation(mod_2824_inner, "mod_2824");
    Operation_IFC mod_2825_inner <- mkFlatten(0);
    Operation_IFC mod_2825 <- mkDebugOperation(mod_2825_inner, "mod_2825");
    Operation_IFC mod_2826_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2826 <- mkDebugOperation(mod_2826_inner, "mod_2826");
    Operation_IFC mod_2827_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2827 <- mkDebugOperation(mod_2827_inner, "mod_2827");
    PMU_IFC mod_2828_bufferize <- mkPMU(2);
    Operation_IFC mod_2828_inner = mod_2828_bufferize.operation;
    Operation_IFC mod_2828 <- mkDebugOperation(mod_2828_inner, "mod_2828");
    rule rule_3605;
        ChannelMessage t;
        t <- mod_2797.get(0);
        mod_2798.put(0, t);
    endrule
    rule rule_3606;
        ChannelMessage t;
        t <- mod_2827.get(0);
        mod_2794.put(1, t);
    endrule
    rule rule_3607;
        ChannelMessage t;
        t <- mod_2796.get(0);
        mod_2826.put(0, t);
    endrule
    rule rule_3608;
        ChannelMessage t;
        t <- mod_2794.get(1);
        mod_2795.put(0, t);
    endrule
    rule rule_3609;
        ChannelMessage t;
        t <- mod_2795.get(0);
        mod_2820.put(0, t);
    endrule
    rule rule_3610;
        ChannelMessage t;
        t <- mod_2816.get(1);
        mod_2815.put(1, t);
    endrule
    rule rule_3611;
        ChannelMessage t;
        t <- mod_2807.get(0);
        mod_2807.put(1, t);
    endrule
    rule rule_3612;
        ChannelMessage t;
        t <- mod_2814.get(0);
        mod_2813.put(0, t);
    endrule
    rule rule_3613;
        ChannelMessage t;
        t <- mod_2819.get(0);
        mod_2818.put(0, t);
    endrule
    rule rule_3614;
        ChannelMessage t;
        t <- mod_2789.get(0);
        mod_2790.put(0, t);
    endrule
    rule rule_3615;
        ChannelMessage t;
        t <- mod_2826.get(0);
        mod_2796.put(1, t);
    endrule
    rule rule_3616;
        ChannelMessage t;
        t <- mod_2822.get(0);
        mod_2823.put(0, t);
    endrule
    rule rule_3617;
        ChannelMessage t;
        t <- mod_2816.get(0);
        mod_2817.put(0, t);
    endrule
    rule rule_3618;
        ChannelMessage t;
        t <- mod_2824.get(0);
        mod_2822.put(0, t);
    endrule
    rule rule_3619;
        ChannelMessage t;
        t <- mod_2809.get(0);
        mod_2808.put(1, t);
    endrule
    rule rule_3620;
        ChannelMessage t;
        t <- mod_2822.get(1);
        mod_2797.put(1, t);
    endrule
    rule rule_3621;
        ChannelMessage t;
        t <- mod_2793.get(3);
        mod_2794.put(0, t);
    endrule
    rule rule_3622;
        ChannelMessage t;
        t <- mod_2796.get(1);
        mod_2797.put(0, t);
    endrule
    rule rule_3623;
        ChannelMessage t;
        t <- mod_2818.get(0);
        mod_2816.put(0, t);
    endrule
    rule rule_3624;
        ChannelMessage t;
        t <- mod_2802.get(0);
        mod_2803.put(0, t);
    endrule
    rule rule_3625;
        ChannelMessage t;
        t <- mod_2804.get(0);
        mod_2806.put(0, t);
    endrule
    rule rule_3626;
        ChannelMessage t;
        t <- mod_2799.get(0);
        mod_2800.put(0, t);
    endrule
    rule rule_3627;
        ChannelMessage t;
        t <- mod_2801.get(0);
        mod_2802.put(0, t);
    endrule
    rule rule_3628;
        ChannelMessage t;
        t <- mod_2800.get(0);
        mod_2812.put(0, t);
    endrule
    rule rule_3629;
        ChannelMessage t;
        t <- mod_2794.get(0);
        mod_2827.put(0, t);
    endrule
    rule rule_3630;
        ChannelMessage t;
        t <- mod_2811.get(0);
        mod_2810.put(0, t);
    endrule
    rule rule_3631;
        ChannelMessage t;
        t <- mod_2820.get(0);
        mod_2821.put(0, t);
    endrule
    rule rule_3632;
        ChannelMessage t;
        t <- mod_2825.get(0);
        mod_2824.put(0, t);
    endrule
    rule rule_3633;
        ChannelMessage t;
        t <- mod_2828.get(1);
        mod_2792.put(1, t);
    endrule
    rule rule_3634;
        ChannelMessage t;
        t <- mod_2823.get(0);
        mod_2822.put(1, t);
    endrule
    rule rule_3635;
        ChannelMessage t;
        t <- mod_2806.get(1);
        mod_2804.put(1, t);
    endrule
    rule rule_3636;
        ChannelMessage t;
        t <- mod_2807.get(1);
        mod_2803.put(1, t);
    endrule
    rule rule_3637;
        ChannelMessage t;
        t <- mod_2800.get(1);
        mod_2801.put(0, t);
    endrule
    rule rule_3638;
        ChannelMessage t;
        t <- mod_2810.get(0);
        mod_2808.put(0, t);
    endrule
    rule rule_3639;
        ChannelMessage t;
        t <- mod_2817.get(0);
        mod_2816.put(1, t);
    endrule
    rule rule_3640;
        ChannelMessage t;
        t <- mod_2803.get(1);
        mod_2804.put(0, t);
    endrule
    rule rule_3641;
        ChannelMessage t;
        t <- mod_2803.get(0);
        mod_2807.put(0, t);
    endrule
    rule rule_3642;
        ChannelMessage t;
        t <- mod_2806.get(0);
        mod_2806.put(1, t);
    endrule
    rule rule_3643;
        ChannelMessage t;
        t <- mod_2795.get(1);
        mod_2796.put(0, t);
    endrule
    rule rule_3644;
        ChannelMessage t;
        t <- mod_2828.get(0);
        mod_2828.put(1, t);
    endrule
    rule rule_3645;
        ChannelMessage t;
        t <- mod_2790.get(0);
        mod_2791.put(0, t);
    endrule
    rule rule_3646;
        ChannelMessage t;
        t <- mod_2791.get(0);
        mod_2792.put(0, t);
    endrule
    rule rule_3647;
        ChannelMessage t;
        t <- mod_2804.get(1);
        mod_2805.put(1, t);
    endrule
    rule rule_3648;
        ChannelMessage t;
        t <- mod_2813.get(0);
        mod_2799.put(1, t);
    endrule
    rule rule_3649;
        ChannelMessage t;
        t <- mod_2808.get(0);
        mod_2809.put(0, t);
    endrule
    rule rule_3650;
        ChannelMessage t;
        t <- mod_2815.get(0);
        mod_2814.put(0, t);
    endrule
    rule rule_3651;
        ChannelMessage t;
        t <- mod_2812.get(0);
        mod_2800.put(1, t);
    endrule
    rule rule_3652;
        ChannelMessage t;
        t <- mod_2792.get(0);
        mod_2828.put(0, t);
    endrule
    rule rule_3653;
        ChannelMessage t;
        t <- mod_2798.get(0);
        mod_2799.put(0, t);
    endrule
    rule rule_3654;
        ChannelMessage t;
        t <- mod_2792.get(1);
        mod_2793.put(0, t);
    endrule
    rule rule_3655;
        ChannelMessage t;
        t <- mod_2820.get(1);
        mod_2815.put(0, t);
    endrule
    rule rule_3656;
        ChannelMessage t;
        t <- mod_2808.get(1);
        mod_2801.put(1, t);
    endrule
    rule rule_3657;
        ChannelMessage t;
        t <- mod_2821.get(0);
        mod_2820.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2789.put(0, t);
        end
        if (i == 1) begin
            mod_2805.put(0, t);
        end
        if (i == 2) begin
            mod_2811.put(0, t);
        end
        if (i == 3) begin
            mod_2819.put(0, t);
        end
        if (i == 4) begin
            mod_2825.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_2793.get(0);
        end
        if (i == 1) begin
            t <- mod_2793.get(1);
        end
        if (i == 2) begin
            t <- mod_2793.get(2);
        end
        if (i == 0) begin
            t <- mod_2805.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6103 (Operation_IFC);
    Operation_IFC mod_2830_inner <- mkReshape(2, 64);
    Operation_IFC mod_2830 <- mkDebugOperation(mod_2830_inner, "mod_2830");
    Operation_IFC mod_2831_inner <- mkFlatten(1);
    Operation_IFC mod_2831 <- mkDebugOperation(mod_2831_inner, "mod_2831");
    Operation_IFC mod_2832_inner <- mkFlatten(2);
    Operation_IFC mod_2832 <- mkDebugOperation(mod_2832_inner, "mod_2832");
    Operation_IFC mod_2833_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2833 <- mkDebugOperation(mod_2833_inner, "mod_2833");
    Broadcast_IFC#(4) mod_2834_inner <- mkBroadcast(4);
    Operation_IFC mod_2834 <- mkDebugOperation(mod_2834_inner.op, "mod_2834");
    PMU_IFC mod_2835_bufferize <- mkPMU(2);
    Operation_IFC mod_2835_inner = mod_2835_bufferize.operation;
    Operation_IFC mod_2835 <- mkDebugOperation(mod_2835_inner, "mod_2835");
    Broadcast_IFC#(2) mod_2836_inner <- mkBroadcast(2);
    Operation_IFC mod_2836 <- mkDebugOperation(mod_2836_inner.op, "mod_2836");
    PMU_IFC mod_2837_bufferize <- mkPMU(1);
    Operation_IFC mod_2837_inner = mod_2837_bufferize.operation;
    Operation_IFC mod_2837 <- mkDebugOperation(mod_2837_inner, "mod_2837");
    Operation_IFC mod_2838_inner <- mkBinaryMap(1087, matmul_t_tile);
    Operation_IFC mod_2838 <- mkDebugOperation(mod_2838_inner, "mod_2838");
    Operation_IFC mod_2839_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2839 <- mkDebugOperation(mod_2839_inner, "mod_2839");
    Operation_IFC mod_2840_inner <- mkBinaryMap(1855, mul_tile);
    Operation_IFC mod_2840 <- mkDebugOperation(mod_2840_inner, "mod_2840");
    PMU_IFC mod_2841_bufferize <- mkPMU(1);
    Operation_IFC mod_2841_inner = mod_2841_bufferize.operation;
    Operation_IFC mod_2841 <- mkDebugOperation(mod_2841_inner, "mod_2841");
    Operation_IFC mod_2842_inner <- mkBinaryMap(2425, matmul_t_tile);
    Operation_IFC mod_2842 <- mkDebugOperation(mod_2842_inner, "mod_2842");
    Operation_IFC mod_2843_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2843 <- mkDebugOperation(mod_2843_inner, "mod_2843");
    Operation_IFC mod_2844_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2844 <- mkDebugOperation(mod_2844_inner, "mod_2844");
    Operation_IFC mod_2845_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2845 <- mkDebugOperation(mod_2845_inner, "mod_2845");
    Operation_IFC mod_2846_inner <- mkBinaryMap(2754, mul_tile);
    Operation_IFC mod_2846 <- mkDebugOperation(mod_2846_inner, "mod_2846");
    PMU_IFC mod_2847_bufferize <- mkPMU(1);
    Operation_IFC mod_2847_inner = mod_2847_bufferize.operation;
    Operation_IFC mod_2847 <- mkDebugOperation(mod_2847_inner, "mod_2847");
    PMU_IFC mod_2848_bufferize <- mkPMU(2);
    Operation_IFC mod_2848_inner = mod_2848_bufferize.operation;
    Operation_IFC mod_2848 <- mkDebugOperation(mod_2848_inner, "mod_2848");
    PMU_IFC mod_2849_bufferize <- mkPMU(2);
    Operation_IFC mod_2849_inner = mod_2849_bufferize.operation;
    Operation_IFC mod_2849 <- mkDebugOperation(mod_2849_inner, "mod_2849");
    Operation_IFC mod_2850_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2850 <- mkDebugOperation(mod_2850_inner, "mod_2850");
    Operation_IFC mod_2851_inner <- mkFlatten(1);
    Operation_IFC mod_2851 <- mkDebugOperation(mod_2851_inner, "mod_2851");
    Operation_IFC mod_2852_inner <- mkFlatten(0);
    Operation_IFC mod_2852 <- mkDebugOperation(mod_2852_inner, "mod_2852");
    Operation_IFC mod_2853_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2853 <- mkDebugOperation(mod_2853_inner, "mod_2853");
    Operation_IFC mod_2854_inner <- mkUnaryMap(1727, silu_tile);
    Operation_IFC mod_2854 <- mkDebugOperation(mod_2854_inner, "mod_2854");
    Operation_IFC mod_2855_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2855 <- mkDebugOperation(mod_2855_inner, "mod_2855");
    Operation_IFC mod_2856_inner <- mkBinaryMap(1599, matmul_t_tile);
    Operation_IFC mod_2856 <- mkDebugOperation(mod_2856_inner, "mod_2856");
    PMU_IFC mod_2857_bufferize <- mkPMU(2);
    Operation_IFC mod_2857_inner = mod_2857_bufferize.operation;
    Operation_IFC mod_2857 <- mkDebugOperation(mod_2857_inner, "mod_2857");
    Operation_IFC mod_2858_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2858 <- mkDebugOperation(mod_2858_inner, "mod_2858");
    Operation_IFC mod_2859_inner <- mkFlatten(1);
    Operation_IFC mod_2859 <- mkDebugOperation(mod_2859_inner, "mod_2859");
    Operation_IFC mod_2860_inner <- mkFlatten(0);
    Operation_IFC mod_2860 <- mkDebugOperation(mod_2860_inner, "mod_2860");
    PMU_IFC mod_2861_bufferize <- mkPMU(1);
    Operation_IFC mod_2861_inner = mod_2861_bufferize.operation;
    Operation_IFC mod_2861 <- mkDebugOperation(mod_2861_inner, "mod_2861");
    Operation_IFC mod_2862_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2862 <- mkDebugOperation(mod_2862_inner, "mod_2862");
    PMU_IFC mod_2863_bufferize <- mkPMU(2);
    Operation_IFC mod_2863_inner = mod_2863_bufferize.operation;
    Operation_IFC mod_2863 <- mkDebugOperation(mod_2863_inner, "mod_2863");
    Operation_IFC mod_2864_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2864 <- mkDebugOperation(mod_2864_inner, "mod_2864");
    Operation_IFC mod_2865_inner <- mkFlatten(1);
    Operation_IFC mod_2865 <- mkDebugOperation(mod_2865_inner, "mod_2865");
    Operation_IFC mod_2866_inner <- mkFlatten(0);
    Operation_IFC mod_2866 <- mkDebugOperation(mod_2866_inner, "mod_2866");
    Operation_IFC mod_2867_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2867 <- mkDebugOperation(mod_2867_inner, "mod_2867");
    Operation_IFC mod_2868_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2868 <- mkDebugOperation(mod_2868_inner, "mod_2868");
    PMU_IFC mod_2869_bufferize <- mkPMU(2);
    Operation_IFC mod_2869_inner = mod_2869_bufferize.operation;
    Operation_IFC mod_2869 <- mkDebugOperation(mod_2869_inner, "mod_2869");
    rule rule_3658;
        ChannelMessage t;
        t <- mod_2833.get(0);
        mod_2869.put(0, t);
    endrule
    rule rule_3659;
        ChannelMessage t;
        t <- mod_2851.get(0);
        mod_2849.put(0, t);
    endrule
    rule rule_3660;
        ChannelMessage t;
        t <- mod_2845.get(0);
        mod_2847.put(0, t);
    endrule
    rule rule_3661;
        ChannelMessage t;
        t <- mod_2863.get(1);
        mod_2838.put(1, t);
    endrule
    rule rule_3662;
        ChannelMessage t;
        t <- mod_2869.get(1);
        mod_2833.put(1, t);
    endrule
    rule rule_3663;
        ChannelMessage t;
        t <- mod_2838.get(0);
        mod_2839.put(0, t);
    endrule
    rule rule_3664;
        ChannelMessage t;
        t <- mod_2836.get(1);
        mod_2837.put(0, t);
    endrule
    rule rule_3665;
        ChannelMessage t;
        t <- mod_2863.get(0);
        mod_2864.put(0, t);
    endrule
    rule rule_3666;
        ChannelMessage t;
        t <- mod_2843.get(0);
        mod_2844.put(0, t);
    endrule
    rule rule_3667;
        ChannelMessage t;
        t <- mod_2844.get(1);
        mod_2845.put(0, t);
    endrule
    rule rule_3668;
        ChannelMessage t;
        t <- mod_2856.get(0);
        mod_2855.put(0, t);
    endrule
    rule rule_3669;
        ChannelMessage t;
        t <- mod_2857.get(0);
        mod_2858.put(0, t);
    endrule
    rule rule_3670;
        ChannelMessage t;
        t <- mod_2837.get(1);
        mod_2838.put(0, t);
    endrule
    rule rule_3671;
        ChannelMessage t;
        t <- mod_2847.get(1);
        mod_2845.put(1, t);
    endrule
    rule rule_3672;
        ChannelMessage t;
        t <- mod_2836.get(0);
        mod_2861.put(0, t);
    endrule
    rule rule_3673;
        ChannelMessage t;
        t <- mod_2867.get(0);
        mod_2837.put(1, t);
    endrule
    rule rule_3674;
        ChannelMessage t;
        t <- mod_2864.get(0);
        mod_2863.put(1, t);
    endrule
    rule rule_3675;
        ChannelMessage t;
        t <- mod_2835.get(0);
        mod_2868.put(0, t);
    endrule
    rule rule_3676;
        ChannelMessage t;
        t <- mod_2860.get(0);
        mod_2859.put(0, t);
    endrule
    rule rule_3677;
        ChannelMessage t;
        t <- mod_2840.get(0);
        mod_2841.put(0, t);
    endrule
    rule rule_3678;
        ChannelMessage t;
        t <- mod_2866.get(0);
        mod_2865.put(0, t);
    endrule
    rule rule_3679;
        ChannelMessage t;
        t <- mod_2861.get(0);
        mod_2862.put(0, t);
    endrule
    rule rule_3680;
        ChannelMessage t;
        t <- mod_2834.get(3);
        mod_2835.put(0, t);
    endrule
    rule rule_3681;
        ChannelMessage t;
        t <- mod_2844.get(0);
        mod_2848.put(0, t);
    endrule
    rule rule_3682;
        ChannelMessage t;
        t <- mod_2848.get(0);
        mod_2848.put(1, t);
    endrule
    rule rule_3683;
        ChannelMessage t;
        t <- mod_2852.get(0);
        mod_2851.put(0, t);
    endrule
    rule rule_3684;
        ChannelMessage t;
        t <- mod_2862.get(0);
        mod_2861.put(1, t);
    endrule
    rule rule_3685;
        ChannelMessage t;
        t <- mod_2858.get(0);
        mod_2857.put(1, t);
    endrule
    rule rule_3686;
        ChannelMessage t;
        t <- mod_2855.get(0);
        mod_2854.put(0, t);
    endrule
    rule rule_3687;
        ChannelMessage t;
        t <- mod_2832.get(0);
        mod_2833.put(0, t);
    endrule
    rule rule_3688;
        ChannelMessage t;
        t <- mod_2859.get(0);
        mod_2857.put(0, t);
    endrule
    rule rule_3689;
        ChannelMessage t;
        t <- mod_2841.get(0);
        mod_2853.put(0, t);
    endrule
    rule rule_3690;
        ChannelMessage t;
        t <- mod_2841.get(1);
        mod_2842.put(0, t);
    endrule
    rule rule_3691;
        ChannelMessage t;
        t <- mod_2837.get(0);
        mod_2867.put(0, t);
    endrule
    rule rule_3692;
        ChannelMessage t;
        t <- mod_2868.get(0);
        mod_2835.put(1, t);
    endrule
    rule rule_3693;
        ChannelMessage t;
        t <- mod_2830.get(0);
        mod_2831.put(0, t);
    endrule
    rule rule_3694;
        ChannelMessage t;
        t <- mod_2849.get(0);
        mod_2850.put(0, t);
    endrule
    rule rule_3695;
        ChannelMessage t;
        t <- mod_2833.get(1);
        mod_2834.put(0, t);
    endrule
    rule rule_3696;
        ChannelMessage t;
        t <- mod_2842.get(0);
        mod_2843.put(0, t);
    endrule
    rule rule_3697;
        ChannelMessage t;
        t <- mod_2857.get(1);
        mod_2856.put(1, t);
    endrule
    rule rule_3698;
        ChannelMessage t;
        t <- mod_2865.get(0);
        mod_2863.put(0, t);
    endrule
    rule rule_3699;
        ChannelMessage t;
        t <- mod_2848.get(1);
        mod_2844.put(1, t);
    endrule
    rule rule_3700;
        ChannelMessage t;
        t <- mod_2831.get(0);
        mod_2832.put(0, t);
    endrule
    rule rule_3701;
        ChannelMessage t;
        t <- mod_2849.get(1);
        mod_2842.put(1, t);
    endrule
    rule rule_3702;
        ChannelMessage t;
        t <- mod_2853.get(0);
        mod_2841.put(1, t);
    endrule
    rule rule_3703;
        ChannelMessage t;
        t <- mod_2854.get(0);
        mod_2840.put(1, t);
    endrule
    rule rule_3704;
        ChannelMessage t;
        t <- mod_2845.get(1);
        mod_2846.put(1, t);
    endrule
    rule rule_3705;
        ChannelMessage t;
        t <- mod_2839.get(0);
        mod_2840.put(0, t);
    endrule
    rule rule_3706;
        ChannelMessage t;
        t <- mod_2835.get(1);
        mod_2836.put(0, t);
    endrule
    rule rule_3707;
        ChannelMessage t;
        t <- mod_2869.get(0);
        mod_2869.put(1, t);
    endrule
    rule rule_3708;
        ChannelMessage t;
        t <- mod_2847.get(0);
        mod_2847.put(1, t);
    endrule
    rule rule_3709;
        ChannelMessage t;
        t <- mod_2850.get(0);
        mod_2849.put(1, t);
    endrule
    rule rule_3710;
        ChannelMessage t;
        t <- mod_2861.get(1);
        mod_2856.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2830.put(0, t);
        end
        if (i == 1) begin
            mod_2846.put(0, t);
        end
        if (i == 2) begin
            mod_2852.put(0, t);
        end
        if (i == 3) begin
            mod_2860.put(0, t);
        end
        if (i == 4) begin
            mod_2866.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_2834.get(0);
        end
        if (i == 2) begin
            t <- mod_2834.get(1);
        end
        if (i == 1) begin
            t <- mod_2834.get(2);
        end
        if (i == 3) begin
            t <- mod_2846.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6104 (Operation_IFC);
    Operation_IFC mod_2871_inner <- mkReshape(2, 64);
    Operation_IFC mod_2871 <- mkDebugOperation(mod_2871_inner, "mod_2871");
    Operation_IFC mod_2872_inner <- mkFlatten(1);
    Operation_IFC mod_2872 <- mkDebugOperation(mod_2872_inner, "mod_2872");
    Operation_IFC mod_2873_inner <- mkFlatten(2);
    Operation_IFC mod_2873 <- mkDebugOperation(mod_2873_inner, "mod_2873");
    Operation_IFC mod_2874_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2874 <- mkDebugOperation(mod_2874_inner, "mod_2874");
    Broadcast_IFC#(4) mod_2875_inner <- mkBroadcast(4);
    Operation_IFC mod_2875 <- mkDebugOperation(mod_2875_inner.op, "mod_2875");
    PMU_IFC mod_2876_bufferize <- mkPMU(2);
    Operation_IFC mod_2876_inner = mod_2876_bufferize.operation;
    Operation_IFC mod_2876 <- mkDebugOperation(mod_2876_inner, "mod_2876");
    Broadcast_IFC#(2) mod_2877_inner <- mkBroadcast(2);
    Operation_IFC mod_2877 <- mkDebugOperation(mod_2877_inner.op, "mod_2877");
    PMU_IFC mod_2878_bufferize <- mkPMU(1);
    Operation_IFC mod_2878_inner = mod_2878_bufferize.operation;
    Operation_IFC mod_2878 <- mkDebugOperation(mod_2878_inner, "mod_2878");
    Operation_IFC mod_2879_inner <- mkBinaryMap(1086, matmul_t_tile);
    Operation_IFC mod_2879 <- mkDebugOperation(mod_2879_inner, "mod_2879");
    Operation_IFC mod_2880_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2880 <- mkDebugOperation(mod_2880_inner, "mod_2880");
    Operation_IFC mod_2881_inner <- mkBinaryMap(1854, mul_tile);
    Operation_IFC mod_2881 <- mkDebugOperation(mod_2881_inner, "mod_2881");
    PMU_IFC mod_2882_bufferize <- mkPMU(1);
    Operation_IFC mod_2882_inner = mod_2882_bufferize.operation;
    Operation_IFC mod_2882 <- mkDebugOperation(mod_2882_inner, "mod_2882");
    Operation_IFC mod_2883_inner <- mkBinaryMap(2423, matmul_t_tile);
    Operation_IFC mod_2883 <- mkDebugOperation(mod_2883_inner, "mod_2883");
    Operation_IFC mod_2884_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2884 <- mkDebugOperation(mod_2884_inner, "mod_2884");
    Operation_IFC mod_2885_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2885 <- mkDebugOperation(mod_2885_inner, "mod_2885");
    Operation_IFC mod_2886_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2886 <- mkDebugOperation(mod_2886_inner, "mod_2886");
    Operation_IFC mod_2887_inner <- mkBinaryMap(2753, mul_tile);
    Operation_IFC mod_2887 <- mkDebugOperation(mod_2887_inner, "mod_2887");
    PMU_IFC mod_2888_bufferize <- mkPMU(1);
    Operation_IFC mod_2888_inner = mod_2888_bufferize.operation;
    Operation_IFC mod_2888 <- mkDebugOperation(mod_2888_inner, "mod_2888");
    PMU_IFC mod_2889_bufferize <- mkPMU(2);
    Operation_IFC mod_2889_inner = mod_2889_bufferize.operation;
    Operation_IFC mod_2889 <- mkDebugOperation(mod_2889_inner, "mod_2889");
    PMU_IFC mod_2890_bufferize <- mkPMU(2);
    Operation_IFC mod_2890_inner = mod_2890_bufferize.operation;
    Operation_IFC mod_2890 <- mkDebugOperation(mod_2890_inner, "mod_2890");
    Operation_IFC mod_2891_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2891 <- mkDebugOperation(mod_2891_inner, "mod_2891");
    Operation_IFC mod_2892_inner <- mkFlatten(1);
    Operation_IFC mod_2892 <- mkDebugOperation(mod_2892_inner, "mod_2892");
    Operation_IFC mod_2893_inner <- mkFlatten(0);
    Operation_IFC mod_2893 <- mkDebugOperation(mod_2893_inner, "mod_2893");
    Operation_IFC mod_2894_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2894 <- mkDebugOperation(mod_2894_inner, "mod_2894");
    Operation_IFC mod_2895_inner <- mkUnaryMap(1726, silu_tile);
    Operation_IFC mod_2895 <- mkDebugOperation(mod_2895_inner, "mod_2895");
    Operation_IFC mod_2896_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2896 <- mkDebugOperation(mod_2896_inner, "mod_2896");
    Operation_IFC mod_2897_inner <- mkBinaryMap(1598, matmul_t_tile);
    Operation_IFC mod_2897 <- mkDebugOperation(mod_2897_inner, "mod_2897");
    PMU_IFC mod_2898_bufferize <- mkPMU(2);
    Operation_IFC mod_2898_inner = mod_2898_bufferize.operation;
    Operation_IFC mod_2898 <- mkDebugOperation(mod_2898_inner, "mod_2898");
    Operation_IFC mod_2899_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2899 <- mkDebugOperation(mod_2899_inner, "mod_2899");
    Operation_IFC mod_2900_inner <- mkFlatten(1);
    Operation_IFC mod_2900 <- mkDebugOperation(mod_2900_inner, "mod_2900");
    Operation_IFC mod_2901_inner <- mkFlatten(0);
    Operation_IFC mod_2901 <- mkDebugOperation(mod_2901_inner, "mod_2901");
    PMU_IFC mod_2902_bufferize <- mkPMU(1);
    Operation_IFC mod_2902_inner = mod_2902_bufferize.operation;
    Operation_IFC mod_2902 <- mkDebugOperation(mod_2902_inner, "mod_2902");
    Operation_IFC mod_2903_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2903 <- mkDebugOperation(mod_2903_inner, "mod_2903");
    PMU_IFC mod_2904_bufferize <- mkPMU(2);
    Operation_IFC mod_2904_inner = mod_2904_bufferize.operation;
    Operation_IFC mod_2904 <- mkDebugOperation(mod_2904_inner, "mod_2904");
    Operation_IFC mod_2905_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2905 <- mkDebugOperation(mod_2905_inner, "mod_2905");
    Operation_IFC mod_2906_inner <- mkFlatten(1);
    Operation_IFC mod_2906 <- mkDebugOperation(mod_2906_inner, "mod_2906");
    Operation_IFC mod_2907_inner <- mkFlatten(0);
    Operation_IFC mod_2907 <- mkDebugOperation(mod_2907_inner, "mod_2907");
    Operation_IFC mod_2908_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2908 <- mkDebugOperation(mod_2908_inner, "mod_2908");
    Operation_IFC mod_2909_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2909 <- mkDebugOperation(mod_2909_inner, "mod_2909");
    PMU_IFC mod_2910_bufferize <- mkPMU(2);
    Operation_IFC mod_2910_inner = mod_2910_bufferize.operation;
    Operation_IFC mod_2910 <- mkDebugOperation(mod_2910_inner, "mod_2910");
    rule rule_3711;
        ChannelMessage t;
        t <- mod_2886.get(0);
        mod_2888.put(0, t);
    endrule
    rule rule_3712;
        ChannelMessage t;
        t <- mod_2877.get(1);
        mod_2878.put(0, t);
    endrule
    rule rule_3713;
        ChannelMessage t;
        t <- mod_2888.get(0);
        mod_2888.put(1, t);
    endrule
    rule rule_3714;
        ChannelMessage t;
        t <- mod_2894.get(0);
        mod_2882.put(1, t);
    endrule
    rule rule_3715;
        ChannelMessage t;
        t <- mod_2904.get(0);
        mod_2905.put(0, t);
    endrule
    rule rule_3716;
        ChannelMessage t;
        t <- mod_2878.get(0);
        mod_2908.put(0, t);
    endrule
    rule rule_3717;
        ChannelMessage t;
        t <- mod_2881.get(0);
        mod_2882.put(0, t);
    endrule
    rule rule_3718;
        ChannelMessage t;
        t <- mod_2885.get(1);
        mod_2886.put(0, t);
    endrule
    rule rule_3719;
        ChannelMessage t;
        t <- mod_2895.get(0);
        mod_2881.put(1, t);
    endrule
    rule rule_3720;
        ChannelMessage t;
        t <- mod_2908.get(0);
        mod_2878.put(1, t);
    endrule
    rule rule_3721;
        ChannelMessage t;
        t <- mod_2885.get(0);
        mod_2889.put(0, t);
    endrule
    rule rule_3722;
        ChannelMessage t;
        t <- mod_2886.get(1);
        mod_2887.put(1, t);
    endrule
    rule rule_3723;
        ChannelMessage t;
        t <- mod_2874.get(0);
        mod_2910.put(0, t);
    endrule
    rule rule_3724;
        ChannelMessage t;
        t <- mod_2879.get(0);
        mod_2880.put(0, t);
    endrule
    rule rule_3725;
        ChannelMessage t;
        t <- mod_2907.get(0);
        mod_2906.put(0, t);
    endrule
    rule rule_3726;
        ChannelMessage t;
        t <- mod_2872.get(0);
        mod_2873.put(0, t);
    endrule
    rule rule_3727;
        ChannelMessage t;
        t <- mod_2889.get(1);
        mod_2885.put(1, t);
    endrule
    rule rule_3728;
        ChannelMessage t;
        t <- mod_2906.get(0);
        mod_2904.put(0, t);
    endrule
    rule rule_3729;
        ChannelMessage t;
        t <- mod_2900.get(0);
        mod_2898.put(0, t);
    endrule
    rule rule_3730;
        ChannelMessage t;
        t <- mod_2904.get(1);
        mod_2879.put(1, t);
    endrule
    rule rule_3731;
        ChannelMessage t;
        t <- mod_2889.get(0);
        mod_2889.put(1, t);
    endrule
    rule rule_3732;
        ChannelMessage t;
        t <- mod_2902.get(1);
        mod_2897.put(0, t);
    endrule
    rule rule_3733;
        ChannelMessage t;
        t <- mod_2892.get(0);
        mod_2890.put(0, t);
    endrule
    rule rule_3734;
        ChannelMessage t;
        t <- mod_2888.get(1);
        mod_2886.put(1, t);
    endrule
    rule rule_3735;
        ChannelMessage t;
        t <- mod_2905.get(0);
        mod_2904.put(1, t);
    endrule
    rule rule_3736;
        ChannelMessage t;
        t <- mod_2876.get(1);
        mod_2877.put(0, t);
    endrule
    rule rule_3737;
        ChannelMessage t;
        t <- mod_2910.get(0);
        mod_2910.put(1, t);
    endrule
    rule rule_3738;
        ChannelMessage t;
        t <- mod_2897.get(0);
        mod_2896.put(0, t);
    endrule
    rule rule_3739;
        ChannelMessage t;
        t <- mod_2896.get(0);
        mod_2895.put(0, t);
    endrule
    rule rule_3740;
        ChannelMessage t;
        t <- mod_2873.get(0);
        mod_2874.put(0, t);
    endrule
    rule rule_3741;
        ChannelMessage t;
        t <- mod_2898.get(0);
        mod_2899.put(0, t);
    endrule
    rule rule_3742;
        ChannelMessage t;
        t <- mod_2874.get(1);
        mod_2875.put(0, t);
    endrule
    rule rule_3743;
        ChannelMessage t;
        t <- mod_2882.get(1);
        mod_2883.put(0, t);
    endrule
    rule rule_3744;
        ChannelMessage t;
        t <- mod_2875.get(3);
        mod_2876.put(0, t);
    endrule
    rule rule_3745;
        ChannelMessage t;
        t <- mod_2880.get(0);
        mod_2881.put(0, t);
    endrule
    rule rule_3746;
        ChannelMessage t;
        t <- mod_2884.get(0);
        mod_2885.put(0, t);
    endrule
    rule rule_3747;
        ChannelMessage t;
        t <- mod_2877.get(0);
        mod_2902.put(0, t);
    endrule
    rule rule_3748;
        ChannelMessage t;
        t <- mod_2876.get(0);
        mod_2909.put(0, t);
    endrule
    rule rule_3749;
        ChannelMessage t;
        t <- mod_2883.get(0);
        mod_2884.put(0, t);
    endrule
    rule rule_3750;
        ChannelMessage t;
        t <- mod_2903.get(0);
        mod_2902.put(1, t);
    endrule
    rule rule_3751;
        ChannelMessage t;
        t <- mod_2882.get(0);
        mod_2894.put(0, t);
    endrule
    rule rule_3752;
        ChannelMessage t;
        t <- mod_2890.get(0);
        mod_2891.put(0, t);
    endrule
    rule rule_3753;
        ChannelMessage t;
        t <- mod_2898.get(1);
        mod_2897.put(1, t);
    endrule
    rule rule_3754;
        ChannelMessage t;
        t <- mod_2878.get(1);
        mod_2879.put(0, t);
    endrule
    rule rule_3755;
        ChannelMessage t;
        t <- mod_2899.get(0);
        mod_2898.put(1, t);
    endrule
    rule rule_3756;
        ChannelMessage t;
        t <- mod_2909.get(0);
        mod_2876.put(1, t);
    endrule
    rule rule_3757;
        ChannelMessage t;
        t <- mod_2871.get(0);
        mod_2872.put(0, t);
    endrule
    rule rule_3758;
        ChannelMessage t;
        t <- mod_2890.get(1);
        mod_2883.put(1, t);
    endrule
    rule rule_3759;
        ChannelMessage t;
        t <- mod_2893.get(0);
        mod_2892.put(0, t);
    endrule
    rule rule_3760;
        ChannelMessage t;
        t <- mod_2901.get(0);
        mod_2900.put(0, t);
    endrule
    rule rule_3761;
        ChannelMessage t;
        t <- mod_2891.get(0);
        mod_2890.put(1, t);
    endrule
    rule rule_3762;
        ChannelMessage t;
        t <- mod_2910.get(1);
        mod_2874.put(1, t);
    endrule
    rule rule_3763;
        ChannelMessage t;
        t <- mod_2902.get(0);
        mod_2903.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2871.put(0, t);
        end
        if (i == 1) begin
            mod_2887.put(0, t);
        end
        if (i == 2) begin
            mod_2893.put(0, t);
        end
        if (i == 3) begin
            mod_2901.put(0, t);
        end
        if (i == 4) begin
            mod_2907.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_2875.get(0);
        end
        if (i == 0) begin
            t <- mod_2875.get(1);
        end
        if (i == 2) begin
            t <- mod_2875.get(2);
        end
        if (i == 1) begin
            t <- mod_2887.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6105 (Operation_IFC);
    Operation_IFC mod_2912_inner <- mkReshape(2, 64);
    Operation_IFC mod_2912 <- mkDebugOperation(mod_2912_inner, "mod_2912");
    Operation_IFC mod_2913_inner <- mkFlatten(1);
    Operation_IFC mod_2913 <- mkDebugOperation(mod_2913_inner, "mod_2913");
    Operation_IFC mod_2914_inner <- mkFlatten(2);
    Operation_IFC mod_2914 <- mkDebugOperation(mod_2914_inner, "mod_2914");
    Operation_IFC mod_2915_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2915 <- mkDebugOperation(mod_2915_inner, "mod_2915");
    Broadcast_IFC#(4) mod_2916_inner <- mkBroadcast(4);
    Operation_IFC mod_2916 <- mkDebugOperation(mod_2916_inner.op, "mod_2916");
    PMU_IFC mod_2917_bufferize <- mkPMU(2);
    Operation_IFC mod_2917_inner = mod_2917_bufferize.operation;
    Operation_IFC mod_2917 <- mkDebugOperation(mod_2917_inner, "mod_2917");
    Broadcast_IFC#(2) mod_2918_inner <- mkBroadcast(2);
    Operation_IFC mod_2918 <- mkDebugOperation(mod_2918_inner.op, "mod_2918");
    PMU_IFC mod_2919_bufferize <- mkPMU(1);
    Operation_IFC mod_2919_inner = mod_2919_bufferize.operation;
    Operation_IFC mod_2919 <- mkDebugOperation(mod_2919_inner, "mod_2919");
    Operation_IFC mod_2920_inner <- mkBinaryMap(1085, matmul_t_tile);
    Operation_IFC mod_2920 <- mkDebugOperation(mod_2920_inner, "mod_2920");
    Operation_IFC mod_2921_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2921 <- mkDebugOperation(mod_2921_inner, "mod_2921");
    Operation_IFC mod_2922_inner <- mkBinaryMap(1853, mul_tile);
    Operation_IFC mod_2922 <- mkDebugOperation(mod_2922_inner, "mod_2922");
    PMU_IFC mod_2923_bufferize <- mkPMU(1);
    Operation_IFC mod_2923_inner = mod_2923_bufferize.operation;
    Operation_IFC mod_2923 <- mkDebugOperation(mod_2923_inner, "mod_2923");
    Operation_IFC mod_2924_inner <- mkBinaryMap(2421, matmul_t_tile);
    Operation_IFC mod_2924 <- mkDebugOperation(mod_2924_inner, "mod_2924");
    Operation_IFC mod_2925_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2925 <- mkDebugOperation(mod_2925_inner, "mod_2925");
    Operation_IFC mod_2926_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2926 <- mkDebugOperation(mod_2926_inner, "mod_2926");
    Operation_IFC mod_2927_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2927 <- mkDebugOperation(mod_2927_inner, "mod_2927");
    Operation_IFC mod_2928_inner <- mkBinaryMap(2752, mul_tile);
    Operation_IFC mod_2928 <- mkDebugOperation(mod_2928_inner, "mod_2928");
    PMU_IFC mod_2929_bufferize <- mkPMU(1);
    Operation_IFC mod_2929_inner = mod_2929_bufferize.operation;
    Operation_IFC mod_2929 <- mkDebugOperation(mod_2929_inner, "mod_2929");
    PMU_IFC mod_2930_bufferize <- mkPMU(2);
    Operation_IFC mod_2930_inner = mod_2930_bufferize.operation;
    Operation_IFC mod_2930 <- mkDebugOperation(mod_2930_inner, "mod_2930");
    PMU_IFC mod_2931_bufferize <- mkPMU(2);
    Operation_IFC mod_2931_inner = mod_2931_bufferize.operation;
    Operation_IFC mod_2931 <- mkDebugOperation(mod_2931_inner, "mod_2931");
    Operation_IFC mod_2932_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2932 <- mkDebugOperation(mod_2932_inner, "mod_2932");
    Operation_IFC mod_2933_inner <- mkFlatten(1);
    Operation_IFC mod_2933 <- mkDebugOperation(mod_2933_inner, "mod_2933");
    Operation_IFC mod_2934_inner <- mkFlatten(0);
    Operation_IFC mod_2934 <- mkDebugOperation(mod_2934_inner, "mod_2934");
    Operation_IFC mod_2935_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2935 <- mkDebugOperation(mod_2935_inner, "mod_2935");
    Operation_IFC mod_2936_inner <- mkUnaryMap(1725, silu_tile);
    Operation_IFC mod_2936 <- mkDebugOperation(mod_2936_inner, "mod_2936");
    Operation_IFC mod_2937_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2937 <- mkDebugOperation(mod_2937_inner, "mod_2937");
    Operation_IFC mod_2938_inner <- mkBinaryMap(1597, matmul_t_tile);
    Operation_IFC mod_2938 <- mkDebugOperation(mod_2938_inner, "mod_2938");
    PMU_IFC mod_2939_bufferize <- mkPMU(2);
    Operation_IFC mod_2939_inner = mod_2939_bufferize.operation;
    Operation_IFC mod_2939 <- mkDebugOperation(mod_2939_inner, "mod_2939");
    Operation_IFC mod_2940_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2940 <- mkDebugOperation(mod_2940_inner, "mod_2940");
    Operation_IFC mod_2941_inner <- mkFlatten(1);
    Operation_IFC mod_2941 <- mkDebugOperation(mod_2941_inner, "mod_2941");
    Operation_IFC mod_2942_inner <- mkFlatten(0);
    Operation_IFC mod_2942 <- mkDebugOperation(mod_2942_inner, "mod_2942");
    PMU_IFC mod_2943_bufferize <- mkPMU(1);
    Operation_IFC mod_2943_inner = mod_2943_bufferize.operation;
    Operation_IFC mod_2943 <- mkDebugOperation(mod_2943_inner, "mod_2943");
    Operation_IFC mod_2944_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2944 <- mkDebugOperation(mod_2944_inner, "mod_2944");
    PMU_IFC mod_2945_bufferize <- mkPMU(2);
    Operation_IFC mod_2945_inner = mod_2945_bufferize.operation;
    Operation_IFC mod_2945 <- mkDebugOperation(mod_2945_inner, "mod_2945");
    Operation_IFC mod_2946_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2946 <- mkDebugOperation(mod_2946_inner, "mod_2946");
    Operation_IFC mod_2947_inner <- mkFlatten(1);
    Operation_IFC mod_2947 <- mkDebugOperation(mod_2947_inner, "mod_2947");
    Operation_IFC mod_2948_inner <- mkFlatten(0);
    Operation_IFC mod_2948 <- mkDebugOperation(mod_2948_inner, "mod_2948");
    Operation_IFC mod_2949_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2949 <- mkDebugOperation(mod_2949_inner, "mod_2949");
    Operation_IFC mod_2950_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2950 <- mkDebugOperation(mod_2950_inner, "mod_2950");
    PMU_IFC mod_2951_bufferize <- mkPMU(2);
    Operation_IFC mod_2951_inner = mod_2951_bufferize.operation;
    Operation_IFC mod_2951 <- mkDebugOperation(mod_2951_inner, "mod_2951");
    rule rule_3764;
        ChannelMessage t;
        t <- mod_2924.get(0);
        mod_2925.put(0, t);
    endrule
    rule rule_3765;
        ChannelMessage t;
        t <- mod_2935.get(0);
        mod_2923.put(1, t);
    endrule
    rule rule_3766;
        ChannelMessage t;
        t <- mod_2944.get(0);
        mod_2943.put(1, t);
    endrule
    rule rule_3767;
        ChannelMessage t;
        t <- mod_2936.get(0);
        mod_2922.put(1, t);
    endrule
    rule rule_3768;
        ChannelMessage t;
        t <- mod_2945.get(1);
        mod_2920.put(1, t);
    endrule
    rule rule_3769;
        ChannelMessage t;
        t <- mod_2927.get(1);
        mod_2928.put(1, t);
    endrule
    rule rule_3770;
        ChannelMessage t;
        t <- mod_2912.get(0);
        mod_2913.put(0, t);
    endrule
    rule rule_3771;
        ChannelMessage t;
        t <- mod_2947.get(0);
        mod_2945.put(0, t);
    endrule
    rule rule_3772;
        ChannelMessage t;
        t <- mod_2938.get(0);
        mod_2937.put(0, t);
    endrule
    rule rule_3773;
        ChannelMessage t;
        t <- mod_2927.get(0);
        mod_2929.put(0, t);
    endrule
    rule rule_3774;
        ChannelMessage t;
        t <- mod_2914.get(0);
        mod_2915.put(0, t);
    endrule
    rule rule_3775;
        ChannelMessage t;
        t <- mod_2919.get(1);
        mod_2920.put(0, t);
    endrule
    rule rule_3776;
        ChannelMessage t;
        t <- mod_2945.get(0);
        mod_2946.put(0, t);
    endrule
    rule rule_3777;
        ChannelMessage t;
        t <- mod_2915.get(0);
        mod_2951.put(0, t);
    endrule
    rule rule_3778;
        ChannelMessage t;
        t <- mod_2941.get(0);
        mod_2939.put(0, t);
    endrule
    rule rule_3779;
        ChannelMessage t;
        t <- mod_2916.get(3);
        mod_2917.put(0, t);
    endrule
    rule rule_3780;
        ChannelMessage t;
        t <- mod_2926.get(0);
        mod_2930.put(0, t);
    endrule
    rule rule_3781;
        ChannelMessage t;
        t <- mod_2917.get(1);
        mod_2918.put(0, t);
    endrule
    rule rule_3782;
        ChannelMessage t;
        t <- mod_2917.get(0);
        mod_2950.put(0, t);
    endrule
    rule rule_3783;
        ChannelMessage t;
        t <- mod_2920.get(0);
        mod_2921.put(0, t);
    endrule
    rule rule_3784;
        ChannelMessage t;
        t <- mod_2937.get(0);
        mod_2936.put(0, t);
    endrule
    rule rule_3785;
        ChannelMessage t;
        t <- mod_2933.get(0);
        mod_2931.put(0, t);
    endrule
    rule rule_3786;
        ChannelMessage t;
        t <- mod_2934.get(0);
        mod_2933.put(0, t);
    endrule
    rule rule_3787;
        ChannelMessage t;
        t <- mod_2919.get(0);
        mod_2949.put(0, t);
    endrule
    rule rule_3788;
        ChannelMessage t;
        t <- mod_2922.get(0);
        mod_2923.put(0, t);
    endrule
    rule rule_3789;
        ChannelMessage t;
        t <- mod_2951.get(1);
        mod_2915.put(1, t);
    endrule
    rule rule_3790;
        ChannelMessage t;
        t <- mod_2931.get(1);
        mod_2924.put(1, t);
    endrule
    rule rule_3791;
        ChannelMessage t;
        t <- mod_2915.get(1);
        mod_2916.put(0, t);
    endrule
    rule rule_3792;
        ChannelMessage t;
        t <- mod_2923.get(1);
        mod_2924.put(0, t);
    endrule
    rule rule_3793;
        ChannelMessage t;
        t <- mod_2930.get(1);
        mod_2926.put(1, t);
    endrule
    rule rule_3794;
        ChannelMessage t;
        t <- mod_2946.get(0);
        mod_2945.put(1, t);
    endrule
    rule rule_3795;
        ChannelMessage t;
        t <- mod_2932.get(0);
        mod_2931.put(1, t);
    endrule
    rule rule_3796;
        ChannelMessage t;
        t <- mod_2918.get(1);
        mod_2919.put(0, t);
    endrule
    rule rule_3797;
        ChannelMessage t;
        t <- mod_2940.get(0);
        mod_2939.put(1, t);
    endrule
    rule rule_3798;
        ChannelMessage t;
        t <- mod_2951.get(0);
        mod_2951.put(1, t);
    endrule
    rule rule_3799;
        ChannelMessage t;
        t <- mod_2926.get(1);
        mod_2927.put(0, t);
    endrule
    rule rule_3800;
        ChannelMessage t;
        t <- mod_2921.get(0);
        mod_2922.put(0, t);
    endrule
    rule rule_3801;
        ChannelMessage t;
        t <- mod_2929.get(0);
        mod_2929.put(1, t);
    endrule
    rule rule_3802;
        ChannelMessage t;
        t <- mod_2930.get(0);
        mod_2930.put(1, t);
    endrule
    rule rule_3803;
        ChannelMessage t;
        t <- mod_2943.get(0);
        mod_2944.put(0, t);
    endrule
    rule rule_3804;
        ChannelMessage t;
        t <- mod_2948.get(0);
        mod_2947.put(0, t);
    endrule
    rule rule_3805;
        ChannelMessage t;
        t <- mod_2943.get(1);
        mod_2938.put(0, t);
    endrule
    rule rule_3806;
        ChannelMessage t;
        t <- mod_2923.get(0);
        mod_2935.put(0, t);
    endrule
    rule rule_3807;
        ChannelMessage t;
        t <- mod_2925.get(0);
        mod_2926.put(0, t);
    endrule
    rule rule_3808;
        ChannelMessage t;
        t <- mod_2949.get(0);
        mod_2919.put(1, t);
    endrule
    rule rule_3809;
        ChannelMessage t;
        t <- mod_2939.get(1);
        mod_2938.put(1, t);
    endrule
    rule rule_3810;
        ChannelMessage t;
        t <- mod_2939.get(0);
        mod_2940.put(0, t);
    endrule
    rule rule_3811;
        ChannelMessage t;
        t <- mod_2918.get(0);
        mod_2943.put(0, t);
    endrule
    rule rule_3812;
        ChannelMessage t;
        t <- mod_2942.get(0);
        mod_2941.put(0, t);
    endrule
    rule rule_3813;
        ChannelMessage t;
        t <- mod_2913.get(0);
        mod_2914.put(0, t);
    endrule
    rule rule_3814;
        ChannelMessage t;
        t <- mod_2929.get(1);
        mod_2927.put(1, t);
    endrule
    rule rule_3815;
        ChannelMessage t;
        t <- mod_2931.get(0);
        mod_2932.put(0, t);
    endrule
    rule rule_3816;
        ChannelMessage t;
        t <- mod_2950.get(0);
        mod_2917.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2912.put(0, t);
        end
        if (i == 1) begin
            mod_2928.put(0, t);
        end
        if (i == 2) begin
            mod_2934.put(0, t);
        end
        if (i == 3) begin
            mod_2942.put(0, t);
        end
        if (i == 4) begin
            mod_2948.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 2) begin
            t <- mod_2916.get(0);
        end
        if (i == 0) begin
            t <- mod_2916.get(1);
        end
        if (i == 1) begin
            t <- mod_2916.get(2);
        end
        if (i == 3) begin
            t <- mod_2928.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6106 (Operation_IFC);
    Operation_IFC mod_2953_inner <- mkReshape(2, 64);
    Operation_IFC mod_2953 <- mkDebugOperation(mod_2953_inner, "mod_2953");
    Operation_IFC mod_2954_inner <- mkFlatten(1);
    Operation_IFC mod_2954 <- mkDebugOperation(mod_2954_inner, "mod_2954");
    Operation_IFC mod_2955_inner <- mkFlatten(2);
    Operation_IFC mod_2955 <- mkDebugOperation(mod_2955_inner, "mod_2955");
    Operation_IFC mod_2956_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2956 <- mkDebugOperation(mod_2956_inner, "mod_2956");
    Broadcast_IFC#(4) mod_2957_inner <- mkBroadcast(4);
    Operation_IFC mod_2957 <- mkDebugOperation(mod_2957_inner.op, "mod_2957");
    PMU_IFC mod_2958_bufferize <- mkPMU(2);
    Operation_IFC mod_2958_inner = mod_2958_bufferize.operation;
    Operation_IFC mod_2958 <- mkDebugOperation(mod_2958_inner, "mod_2958");
    Broadcast_IFC#(2) mod_2959_inner <- mkBroadcast(2);
    Operation_IFC mod_2959 <- mkDebugOperation(mod_2959_inner.op, "mod_2959");
    PMU_IFC mod_2960_bufferize <- mkPMU(1);
    Operation_IFC mod_2960_inner = mod_2960_bufferize.operation;
    Operation_IFC mod_2960 <- mkDebugOperation(mod_2960_inner, "mod_2960");
    Operation_IFC mod_2961_inner <- mkBinaryMap(1084, matmul_t_tile);
    Operation_IFC mod_2961 <- mkDebugOperation(mod_2961_inner, "mod_2961");
    Operation_IFC mod_2962_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2962 <- mkDebugOperation(mod_2962_inner, "mod_2962");
    Operation_IFC mod_2963_inner <- mkBinaryMap(1852, mul_tile);
    Operation_IFC mod_2963 <- mkDebugOperation(mod_2963_inner, "mod_2963");
    PMU_IFC mod_2964_bufferize <- mkPMU(1);
    Operation_IFC mod_2964_inner = mod_2964_bufferize.operation;
    Operation_IFC mod_2964 <- mkDebugOperation(mod_2964_inner, "mod_2964");
    Operation_IFC mod_2965_inner <- mkBinaryMap(2419, matmul_t_tile);
    Operation_IFC mod_2965 <- mkDebugOperation(mod_2965_inner, "mod_2965");
    Operation_IFC mod_2966_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2966 <- mkDebugOperation(mod_2966_inner, "mod_2966");
    Operation_IFC mod_2967_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_2967 <- mkDebugOperation(mod_2967_inner, "mod_2967");
    Operation_IFC mod_2968_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_2968 <- mkDebugOperation(mod_2968_inner, "mod_2968");
    Operation_IFC mod_2969_inner <- mkBinaryMap(2751, mul_tile);
    Operation_IFC mod_2969 <- mkDebugOperation(mod_2969_inner, "mod_2969");
    PMU_IFC mod_2970_bufferize <- mkPMU(1);
    Operation_IFC mod_2970_inner = mod_2970_bufferize.operation;
    Operation_IFC mod_2970 <- mkDebugOperation(mod_2970_inner, "mod_2970");
    PMU_IFC mod_2971_bufferize <- mkPMU(2);
    Operation_IFC mod_2971_inner = mod_2971_bufferize.operation;
    Operation_IFC mod_2971 <- mkDebugOperation(mod_2971_inner, "mod_2971");
    PMU_IFC mod_2972_bufferize <- mkPMU(2);
    Operation_IFC mod_2972_inner = mod_2972_bufferize.operation;
    Operation_IFC mod_2972 <- mkDebugOperation(mod_2972_inner, "mod_2972");
    Operation_IFC mod_2973_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2973 <- mkDebugOperation(mod_2973_inner, "mod_2973");
    Operation_IFC mod_2974_inner <- mkFlatten(1);
    Operation_IFC mod_2974 <- mkDebugOperation(mod_2974_inner, "mod_2974");
    Operation_IFC mod_2975_inner <- mkFlatten(0);
    Operation_IFC mod_2975 <- mkDebugOperation(mod_2975_inner, "mod_2975");
    Operation_IFC mod_2976_inner <- mkRepeatStatic(3);
    Operation_IFC mod_2976 <- mkDebugOperation(mod_2976_inner, "mod_2976");
    Operation_IFC mod_2977_inner <- mkUnaryMap(1724, silu_tile);
    Operation_IFC mod_2977 <- mkDebugOperation(mod_2977_inner, "mod_2977");
    Operation_IFC mod_2978_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_2978 <- mkDebugOperation(mod_2978_inner, "mod_2978");
    Operation_IFC mod_2979_inner <- mkBinaryMap(1596, matmul_t_tile);
    Operation_IFC mod_2979 <- mkDebugOperation(mod_2979_inner, "mod_2979");
    PMU_IFC mod_2980_bufferize <- mkPMU(2);
    Operation_IFC mod_2980_inner = mod_2980_bufferize.operation;
    Operation_IFC mod_2980 <- mkDebugOperation(mod_2980_inner, "mod_2980");
    Operation_IFC mod_2981_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2981 <- mkDebugOperation(mod_2981_inner, "mod_2981");
    Operation_IFC mod_2982_inner <- mkFlatten(1);
    Operation_IFC mod_2982 <- mkDebugOperation(mod_2982_inner, "mod_2982");
    Operation_IFC mod_2983_inner <- mkFlatten(0);
    Operation_IFC mod_2983 <- mkDebugOperation(mod_2983_inner, "mod_2983");
    PMU_IFC mod_2984_bufferize <- mkPMU(1);
    Operation_IFC mod_2984_inner = mod_2984_bufferize.operation;
    Operation_IFC mod_2984 <- mkDebugOperation(mod_2984_inner, "mod_2984");
    Operation_IFC mod_2985_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2985 <- mkDebugOperation(mod_2985_inner, "mod_2985");
    PMU_IFC mod_2986_bufferize <- mkPMU(2);
    Operation_IFC mod_2986_inner = mod_2986_bufferize.operation;
    Operation_IFC mod_2986 <- mkDebugOperation(mod_2986_inner, "mod_2986");
    Operation_IFC mod_2987_inner <- mkRepeatStatic(8);
    Operation_IFC mod_2987 <- mkDebugOperation(mod_2987_inner, "mod_2987");
    Operation_IFC mod_2988_inner <- mkFlatten(1);
    Operation_IFC mod_2988 <- mkDebugOperation(mod_2988_inner, "mod_2988");
    Operation_IFC mod_2989_inner <- mkFlatten(0);
    Operation_IFC mod_2989 <- mkDebugOperation(mod_2989_inner, "mod_2989");
    Operation_IFC mod_2990_inner <- mkRepeatStatic(16);
    Operation_IFC mod_2990 <- mkDebugOperation(mod_2990_inner, "mod_2990");
    Operation_IFC mod_2991_inner <- mkRepeatStatic(2);
    Operation_IFC mod_2991 <- mkDebugOperation(mod_2991_inner, "mod_2991");
    PMU_IFC mod_2992_bufferize <- mkPMU(2);
    Operation_IFC mod_2992_inner = mod_2992_bufferize.operation;
    Operation_IFC mod_2992 <- mkDebugOperation(mod_2992_inner, "mod_2992");
    rule rule_3817;
        ChannelMessage t;
        t <- mod_2960.get(1);
        mod_2961.put(0, t);
    endrule
    rule rule_3818;
        ChannelMessage t;
        t <- mod_2959.get(0);
        mod_2984.put(0, t);
    endrule
    rule rule_3819;
        ChannelMessage t;
        t <- mod_2955.get(0);
        mod_2956.put(0, t);
    endrule
    rule rule_3820;
        ChannelMessage t;
        t <- mod_2975.get(0);
        mod_2974.put(0, t);
    endrule
    rule rule_3821;
        ChannelMessage t;
        t <- mod_2976.get(0);
        mod_2964.put(1, t);
    endrule
    rule rule_3822;
        ChannelMessage t;
        t <- mod_2988.get(0);
        mod_2986.put(0, t);
    endrule
    rule rule_3823;
        ChannelMessage t;
        t <- mod_2970.get(0);
        mod_2970.put(1, t);
    endrule
    rule rule_3824;
        ChannelMessage t;
        t <- mod_2965.get(0);
        mod_2966.put(0, t);
    endrule
    rule rule_3825;
        ChannelMessage t;
        t <- mod_2956.get(0);
        mod_2992.put(0, t);
    endrule
    rule rule_3826;
        ChannelMessage t;
        t <- mod_2960.get(0);
        mod_2990.put(0, t);
    endrule
    rule rule_3827;
        ChannelMessage t;
        t <- mod_2977.get(0);
        mod_2963.put(1, t);
    endrule
    rule rule_3828;
        ChannelMessage t;
        t <- mod_2986.get(1);
        mod_2961.put(1, t);
    endrule
    rule rule_3829;
        ChannelMessage t;
        t <- mod_2972.get(1);
        mod_2965.put(1, t);
    endrule
    rule rule_3830;
        ChannelMessage t;
        t <- mod_2992.get(0);
        mod_2992.put(1, t);
    endrule
    rule rule_3831;
        ChannelMessage t;
        t <- mod_2974.get(0);
        mod_2972.put(0, t);
    endrule
    rule rule_3832;
        ChannelMessage t;
        t <- mod_2972.get(0);
        mod_2973.put(0, t);
    endrule
    rule rule_3833;
        ChannelMessage t;
        t <- mod_2967.get(1);
        mod_2968.put(0, t);
    endrule
    rule rule_3834;
        ChannelMessage t;
        t <- mod_2971.get(1);
        mod_2967.put(1, t);
    endrule
    rule rule_3835;
        ChannelMessage t;
        t <- mod_2973.get(0);
        mod_2972.put(1, t);
    endrule
    rule rule_3836;
        ChannelMessage t;
        t <- mod_2953.get(0);
        mod_2954.put(0, t);
    endrule
    rule rule_3837;
        ChannelMessage t;
        t <- mod_2992.get(1);
        mod_2956.put(1, t);
    endrule
    rule rule_3838;
        ChannelMessage t;
        t <- mod_2991.get(0);
        mod_2958.put(1, t);
    endrule
    rule rule_3839;
        ChannelMessage t;
        t <- mod_2986.get(0);
        mod_2987.put(0, t);
    endrule
    rule rule_3840;
        ChannelMessage t;
        t <- mod_2958.get(1);
        mod_2959.put(0, t);
    endrule
    rule rule_3841;
        ChannelMessage t;
        t <- mod_2956.get(1);
        mod_2957.put(0, t);
    endrule
    rule rule_3842;
        ChannelMessage t;
        t <- mod_2964.get(1);
        mod_2965.put(0, t);
    endrule
    rule rule_3843;
        ChannelMessage t;
        t <- mod_2957.get(3);
        mod_2958.put(0, t);
    endrule
    rule rule_3844;
        ChannelMessage t;
        t <- mod_2985.get(0);
        mod_2984.put(1, t);
    endrule
    rule rule_3845;
        ChannelMessage t;
        t <- mod_2980.get(1);
        mod_2979.put(1, t);
    endrule
    rule rule_3846;
        ChannelMessage t;
        t <- mod_2979.get(0);
        mod_2978.put(0, t);
    endrule
    rule rule_3847;
        ChannelMessage t;
        t <- mod_2990.get(0);
        mod_2960.put(1, t);
    endrule
    rule rule_3848;
        ChannelMessage t;
        t <- mod_2981.get(0);
        mod_2980.put(1, t);
    endrule
    rule rule_3849;
        ChannelMessage t;
        t <- mod_2964.get(0);
        mod_2976.put(0, t);
    endrule
    rule rule_3850;
        ChannelMessage t;
        t <- mod_2968.get(1);
        mod_2969.put(1, t);
    endrule
    rule rule_3851;
        ChannelMessage t;
        t <- mod_2966.get(0);
        mod_2967.put(0, t);
    endrule
    rule rule_3852;
        ChannelMessage t;
        t <- mod_2959.get(1);
        mod_2960.put(0, t);
    endrule
    rule rule_3853;
        ChannelMessage t;
        t <- mod_2961.get(0);
        mod_2962.put(0, t);
    endrule
    rule rule_3854;
        ChannelMessage t;
        t <- mod_2984.get(0);
        mod_2985.put(0, t);
    endrule
    rule rule_3855;
        ChannelMessage t;
        t <- mod_2967.get(0);
        mod_2971.put(0, t);
    endrule
    rule rule_3856;
        ChannelMessage t;
        t <- mod_2978.get(0);
        mod_2977.put(0, t);
    endrule
    rule rule_3857;
        ChannelMessage t;
        t <- mod_2980.get(0);
        mod_2981.put(0, t);
    endrule
    rule rule_3858;
        ChannelMessage t;
        t <- mod_2989.get(0);
        mod_2988.put(0, t);
    endrule
    rule rule_3859;
        ChannelMessage t;
        t <- mod_2962.get(0);
        mod_2963.put(0, t);
    endrule
    rule rule_3860;
        ChannelMessage t;
        t <- mod_2982.get(0);
        mod_2980.put(0, t);
    endrule
    rule rule_3861;
        ChannelMessage t;
        t <- mod_2984.get(1);
        mod_2979.put(0, t);
    endrule
    rule rule_3862;
        ChannelMessage t;
        t <- mod_2958.get(0);
        mod_2991.put(0, t);
    endrule
    rule rule_3863;
        ChannelMessage t;
        t <- mod_2963.get(0);
        mod_2964.put(0, t);
    endrule
    rule rule_3864;
        ChannelMessage t;
        t <- mod_2954.get(0);
        mod_2955.put(0, t);
    endrule
    rule rule_3865;
        ChannelMessage t;
        t <- mod_2987.get(0);
        mod_2986.put(1, t);
    endrule
    rule rule_3866;
        ChannelMessage t;
        t <- mod_2970.get(1);
        mod_2968.put(1, t);
    endrule
    rule rule_3867;
        ChannelMessage t;
        t <- mod_2983.get(0);
        mod_2982.put(0, t);
    endrule
    rule rule_3868;
        ChannelMessage t;
        t <- mod_2968.get(0);
        mod_2970.put(0, t);
    endrule
    rule rule_3869;
        ChannelMessage t;
        t <- mod_2971.get(0);
        mod_2971.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2953.put(0, t);
        end
        if (i == 1) begin
            mod_2969.put(0, t);
        end
        if (i == 2) begin
            mod_2975.put(0, t);
        end
        if (i == 3) begin
            mod_2983.put(0, t);
        end
        if (i == 4) begin
            mod_2989.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_2957.get(0);
        end
        if (i == 1) begin
            t <- mod_2957.get(1);
        end
        if (i == 2) begin
            t <- mod_2957.get(2);
        end
        if (i == 3) begin
            t <- mod_2969.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6107 (Operation_IFC);
    Operation_IFC mod_2994_inner <- mkReshape(2, 64);
    Operation_IFC mod_2994 <- mkDebugOperation(mod_2994_inner, "mod_2994");
    Operation_IFC mod_2995_inner <- mkFlatten(1);
    Operation_IFC mod_2995 <- mkDebugOperation(mod_2995_inner, "mod_2995");
    Operation_IFC mod_2996_inner <- mkFlatten(2);
    Operation_IFC mod_2996 <- mkDebugOperation(mod_2996_inner, "mod_2996");
    Operation_IFC mod_2997_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_2997 <- mkDebugOperation(mod_2997_inner, "mod_2997");
    Broadcast_IFC#(4) mod_2998_inner <- mkBroadcast(4);
    Operation_IFC mod_2998 <- mkDebugOperation(mod_2998_inner.op, "mod_2998");
    PMU_IFC mod_2999_bufferize <- mkPMU(2);
    Operation_IFC mod_2999_inner = mod_2999_bufferize.operation;
    Operation_IFC mod_2999 <- mkDebugOperation(mod_2999_inner, "mod_2999");
    Broadcast_IFC#(2) mod_3000_inner <- mkBroadcast(2);
    Operation_IFC mod_3000 <- mkDebugOperation(mod_3000_inner.op, "mod_3000");
    PMU_IFC mod_3001_bufferize <- mkPMU(1);
    Operation_IFC mod_3001_inner = mod_3001_bufferize.operation;
    Operation_IFC mod_3001 <- mkDebugOperation(mod_3001_inner, "mod_3001");
    Operation_IFC mod_3002_inner <- mkBinaryMap(1083, matmul_t_tile);
    Operation_IFC mod_3002 <- mkDebugOperation(mod_3002_inner, "mod_3002");
    Operation_IFC mod_3003_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3003 <- mkDebugOperation(mod_3003_inner, "mod_3003");
    Operation_IFC mod_3004_inner <- mkBinaryMap(1851, mul_tile);
    Operation_IFC mod_3004 <- mkDebugOperation(mod_3004_inner, "mod_3004");
    PMU_IFC mod_3005_bufferize <- mkPMU(1);
    Operation_IFC mod_3005_inner = mod_3005_bufferize.operation;
    Operation_IFC mod_3005 <- mkDebugOperation(mod_3005_inner, "mod_3005");
    Operation_IFC mod_3006_inner <- mkBinaryMap(2417, matmul_t_tile);
    Operation_IFC mod_3006 <- mkDebugOperation(mod_3006_inner, "mod_3006");
    Operation_IFC mod_3007_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3007 <- mkDebugOperation(mod_3007_inner, "mod_3007");
    Operation_IFC mod_3008_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3008 <- mkDebugOperation(mod_3008_inner, "mod_3008");
    Operation_IFC mod_3009_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3009 <- mkDebugOperation(mod_3009_inner, "mod_3009");
    Operation_IFC mod_3010_inner <- mkBinaryMap(2750, mul_tile);
    Operation_IFC mod_3010 <- mkDebugOperation(mod_3010_inner, "mod_3010");
    PMU_IFC mod_3011_bufferize <- mkPMU(1);
    Operation_IFC mod_3011_inner = mod_3011_bufferize.operation;
    Operation_IFC mod_3011 <- mkDebugOperation(mod_3011_inner, "mod_3011");
    PMU_IFC mod_3012_bufferize <- mkPMU(2);
    Operation_IFC mod_3012_inner = mod_3012_bufferize.operation;
    Operation_IFC mod_3012 <- mkDebugOperation(mod_3012_inner, "mod_3012");
    PMU_IFC mod_3013_bufferize <- mkPMU(2);
    Operation_IFC mod_3013_inner = mod_3013_bufferize.operation;
    Operation_IFC mod_3013 <- mkDebugOperation(mod_3013_inner, "mod_3013");
    Operation_IFC mod_3014_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3014 <- mkDebugOperation(mod_3014_inner, "mod_3014");
    Operation_IFC mod_3015_inner <- mkFlatten(1);
    Operation_IFC mod_3015 <- mkDebugOperation(mod_3015_inner, "mod_3015");
    Operation_IFC mod_3016_inner <- mkFlatten(0);
    Operation_IFC mod_3016 <- mkDebugOperation(mod_3016_inner, "mod_3016");
    Operation_IFC mod_3017_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3017 <- mkDebugOperation(mod_3017_inner, "mod_3017");
    Operation_IFC mod_3018_inner <- mkUnaryMap(1723, silu_tile);
    Operation_IFC mod_3018 <- mkDebugOperation(mod_3018_inner, "mod_3018");
    Operation_IFC mod_3019_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3019 <- mkDebugOperation(mod_3019_inner, "mod_3019");
    Operation_IFC mod_3020_inner <- mkBinaryMap(1595, matmul_t_tile);
    Operation_IFC mod_3020 <- mkDebugOperation(mod_3020_inner, "mod_3020");
    PMU_IFC mod_3021_bufferize <- mkPMU(2);
    Operation_IFC mod_3021_inner = mod_3021_bufferize.operation;
    Operation_IFC mod_3021 <- mkDebugOperation(mod_3021_inner, "mod_3021");
    Operation_IFC mod_3022_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3022 <- mkDebugOperation(mod_3022_inner, "mod_3022");
    Operation_IFC mod_3023_inner <- mkFlatten(1);
    Operation_IFC mod_3023 <- mkDebugOperation(mod_3023_inner, "mod_3023");
    Operation_IFC mod_3024_inner <- mkFlatten(0);
    Operation_IFC mod_3024 <- mkDebugOperation(mod_3024_inner, "mod_3024");
    PMU_IFC mod_3025_bufferize <- mkPMU(1);
    Operation_IFC mod_3025_inner = mod_3025_bufferize.operation;
    Operation_IFC mod_3025 <- mkDebugOperation(mod_3025_inner, "mod_3025");
    Operation_IFC mod_3026_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3026 <- mkDebugOperation(mod_3026_inner, "mod_3026");
    PMU_IFC mod_3027_bufferize <- mkPMU(2);
    Operation_IFC mod_3027_inner = mod_3027_bufferize.operation;
    Operation_IFC mod_3027 <- mkDebugOperation(mod_3027_inner, "mod_3027");
    Operation_IFC mod_3028_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3028 <- mkDebugOperation(mod_3028_inner, "mod_3028");
    Operation_IFC mod_3029_inner <- mkFlatten(1);
    Operation_IFC mod_3029 <- mkDebugOperation(mod_3029_inner, "mod_3029");
    Operation_IFC mod_3030_inner <- mkFlatten(0);
    Operation_IFC mod_3030 <- mkDebugOperation(mod_3030_inner, "mod_3030");
    Operation_IFC mod_3031_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3031 <- mkDebugOperation(mod_3031_inner, "mod_3031");
    Operation_IFC mod_3032_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3032 <- mkDebugOperation(mod_3032_inner, "mod_3032");
    PMU_IFC mod_3033_bufferize <- mkPMU(2);
    Operation_IFC mod_3033_inner = mod_3033_bufferize.operation;
    Operation_IFC mod_3033 <- mkDebugOperation(mod_3033_inner, "mod_3033");
    rule rule_3870;
        ChannelMessage t;
        t <- mod_3018.get(0);
        mod_3004.put(1, t);
    endrule
    rule rule_3871;
        ChannelMessage t;
        t <- mod_2999.get(1);
        mod_3000.put(0, t);
    endrule
    rule rule_3872;
        ChannelMessage t;
        t <- mod_3011.get(0);
        mod_3011.put(1, t);
    endrule
    rule rule_3873;
        ChannelMessage t;
        t <- mod_3027.get(0);
        mod_3028.put(0, t);
    endrule
    rule rule_3874;
        ChannelMessage t;
        t <- mod_3021.get(1);
        mod_3020.put(1, t);
    endrule
    rule rule_3875;
        ChannelMessage t;
        t <- mod_2999.get(0);
        mod_3032.put(0, t);
    endrule
    rule rule_3876;
        ChannelMessage t;
        t <- mod_3030.get(0);
        mod_3029.put(0, t);
    endrule
    rule rule_3877;
        ChannelMessage t;
        t <- mod_3033.get(1);
        mod_2997.put(1, t);
    endrule
    rule rule_3878;
        ChannelMessage t;
        t <- mod_3015.get(0);
        mod_3013.put(0, t);
    endrule
    rule rule_3879;
        ChannelMessage t;
        t <- mod_3020.get(0);
        mod_3019.put(0, t);
    endrule
    rule rule_3880;
        ChannelMessage t;
        t <- mod_3025.get(1);
        mod_3020.put(0, t);
    endrule
    rule rule_3881;
        ChannelMessage t;
        t <- mod_3001.get(1);
        mod_3002.put(0, t);
    endrule
    rule rule_3882;
        ChannelMessage t;
        t <- mod_2994.get(0);
        mod_2995.put(0, t);
    endrule
    rule rule_3883;
        ChannelMessage t;
        t <- mod_3014.get(0);
        mod_3013.put(1, t);
    endrule
    rule rule_3884;
        ChannelMessage t;
        t <- mod_3013.get(0);
        mod_3014.put(0, t);
    endrule
    rule rule_3885;
        ChannelMessage t;
        t <- mod_3027.get(1);
        mod_3002.put(1, t);
    endrule
    rule rule_3886;
        ChannelMessage t;
        t <- mod_3012.get(0);
        mod_3012.put(1, t);
    endrule
    rule rule_3887;
        ChannelMessage t;
        t <- mod_3008.get(0);
        mod_3012.put(0, t);
    endrule
    rule rule_3888;
        ChannelMessage t;
        t <- mod_3009.get(1);
        mod_3010.put(1, t);
    endrule
    rule rule_3889;
        ChannelMessage t;
        t <- mod_3003.get(0);
        mod_3004.put(0, t);
    endrule
    rule rule_3890;
        ChannelMessage t;
        t <- mod_3022.get(0);
        mod_3021.put(1, t);
    endrule
    rule rule_3891;
        ChannelMessage t;
        t <- mod_3028.get(0);
        mod_3027.put(1, t);
    endrule
    rule rule_3892;
        ChannelMessage t;
        t <- mod_3002.get(0);
        mod_3003.put(0, t);
    endrule
    rule rule_3893;
        ChannelMessage t;
        t <- mod_3031.get(0);
        mod_3001.put(1, t);
    endrule
    rule rule_3894;
        ChannelMessage t;
        t <- mod_3017.get(0);
        mod_3005.put(1, t);
    endrule
    rule rule_3895;
        ChannelMessage t;
        t <- mod_3001.get(0);
        mod_3031.put(0, t);
    endrule
    rule rule_3896;
        ChannelMessage t;
        t <- mod_3011.get(1);
        mod_3009.put(1, t);
    endrule
    rule rule_3897;
        ChannelMessage t;
        t <- mod_3006.get(0);
        mod_3007.put(0, t);
    endrule
    rule rule_3898;
        ChannelMessage t;
        t <- mod_2998.get(3);
        mod_2999.put(0, t);
    endrule
    rule rule_3899;
        ChannelMessage t;
        t <- mod_3024.get(0);
        mod_3023.put(0, t);
    endrule
    rule rule_3900;
        ChannelMessage t;
        t <- mod_3013.get(1);
        mod_3006.put(1, t);
    endrule
    rule rule_3901;
        ChannelMessage t;
        t <- mod_3029.get(0);
        mod_3027.put(0, t);
    endrule
    rule rule_3902;
        ChannelMessage t;
        t <- mod_3016.get(0);
        mod_3015.put(0, t);
    endrule
    rule rule_3903;
        ChannelMessage t;
        t <- mod_3004.get(0);
        mod_3005.put(0, t);
    endrule
    rule rule_3904;
        ChannelMessage t;
        t <- mod_2995.get(0);
        mod_2996.put(0, t);
    endrule
    rule rule_3905;
        ChannelMessage t;
        t <- mod_3021.get(0);
        mod_3022.put(0, t);
    endrule
    rule rule_3906;
        ChannelMessage t;
        t <- mod_3000.get(1);
        mod_3001.put(0, t);
    endrule
    rule rule_3907;
        ChannelMessage t;
        t <- mod_3009.get(0);
        mod_3011.put(0, t);
    endrule
    rule rule_3908;
        ChannelMessage t;
        t <- mod_3025.get(0);
        mod_3026.put(0, t);
    endrule
    rule rule_3909;
        ChannelMessage t;
        t <- mod_3019.get(0);
        mod_3018.put(0, t);
    endrule
    rule rule_3910;
        ChannelMessage t;
        t <- mod_2997.get(0);
        mod_3033.put(0, t);
    endrule
    rule rule_3911;
        ChannelMessage t;
        t <- mod_3007.get(0);
        mod_3008.put(0, t);
    endrule
    rule rule_3912;
        ChannelMessage t;
        t <- mod_2997.get(1);
        mod_2998.put(0, t);
    endrule
    rule rule_3913;
        ChannelMessage t;
        t <- mod_3023.get(0);
        mod_3021.put(0, t);
    endrule
    rule rule_3914;
        ChannelMessage t;
        t <- mod_3005.get(0);
        mod_3017.put(0, t);
    endrule
    rule rule_3915;
        ChannelMessage t;
        t <- mod_3012.get(1);
        mod_3008.put(1, t);
    endrule
    rule rule_3916;
        ChannelMessage t;
        t <- mod_2996.get(0);
        mod_2997.put(0, t);
    endrule
    rule rule_3917;
        ChannelMessage t;
        t <- mod_3005.get(1);
        mod_3006.put(0, t);
    endrule
    rule rule_3918;
        ChannelMessage t;
        t <- mod_3008.get(1);
        mod_3009.put(0, t);
    endrule
    rule rule_3919;
        ChannelMessage t;
        t <- mod_3026.get(0);
        mod_3025.put(1, t);
    endrule
    rule rule_3920;
        ChannelMessage t;
        t <- mod_3000.get(0);
        mod_3025.put(0, t);
    endrule
    rule rule_3921;
        ChannelMessage t;
        t <- mod_3032.get(0);
        mod_2999.put(1, t);
    endrule
    rule rule_3922;
        ChannelMessage t;
        t <- mod_3033.get(0);
        mod_3033.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_2994.put(0, t);
        end
        if (i == 1) begin
            mod_3010.put(0, t);
        end
        if (i == 2) begin
            mod_3016.put(0, t);
        end
        if (i == 3) begin
            mod_3024.put(0, t);
        end
        if (i == 4) begin
            mod_3030.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 2) begin
            t <- mod_2998.get(0);
        end
        if (i == 3) begin
            t <- mod_2998.get(1);
        end
        if (i == 0) begin
            t <- mod_2998.get(2);
        end
        if (i == 1) begin
            t <- mod_3010.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6108 (Operation_IFC);
    Operation_IFC mod_3035_inner <- mkReshape(2, 64);
    Operation_IFC mod_3035 <- mkDebugOperation(mod_3035_inner, "mod_3035");
    Operation_IFC mod_3036_inner <- mkFlatten(1);
    Operation_IFC mod_3036 <- mkDebugOperation(mod_3036_inner, "mod_3036");
    Operation_IFC mod_3037_inner <- mkFlatten(2);
    Operation_IFC mod_3037 <- mkDebugOperation(mod_3037_inner, "mod_3037");
    Operation_IFC mod_3038_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3038 <- mkDebugOperation(mod_3038_inner, "mod_3038");
    Broadcast_IFC#(4) mod_3039_inner <- mkBroadcast(4);
    Operation_IFC mod_3039 <- mkDebugOperation(mod_3039_inner.op, "mod_3039");
    PMU_IFC mod_3040_bufferize <- mkPMU(2);
    Operation_IFC mod_3040_inner = mod_3040_bufferize.operation;
    Operation_IFC mod_3040 <- mkDebugOperation(mod_3040_inner, "mod_3040");
    Broadcast_IFC#(2) mod_3041_inner <- mkBroadcast(2);
    Operation_IFC mod_3041 <- mkDebugOperation(mod_3041_inner.op, "mod_3041");
    PMU_IFC mod_3042_bufferize <- mkPMU(1);
    Operation_IFC mod_3042_inner = mod_3042_bufferize.operation;
    Operation_IFC mod_3042 <- mkDebugOperation(mod_3042_inner, "mod_3042");
    Operation_IFC mod_3043_inner <- mkBinaryMap(1082, matmul_t_tile);
    Operation_IFC mod_3043 <- mkDebugOperation(mod_3043_inner, "mod_3043");
    Operation_IFC mod_3044_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3044 <- mkDebugOperation(mod_3044_inner, "mod_3044");
    Operation_IFC mod_3045_inner <- mkBinaryMap(1850, mul_tile);
    Operation_IFC mod_3045 <- mkDebugOperation(mod_3045_inner, "mod_3045");
    PMU_IFC mod_3046_bufferize <- mkPMU(1);
    Operation_IFC mod_3046_inner = mod_3046_bufferize.operation;
    Operation_IFC mod_3046 <- mkDebugOperation(mod_3046_inner, "mod_3046");
    Operation_IFC mod_3047_inner <- mkBinaryMap(2415, matmul_t_tile);
    Operation_IFC mod_3047 <- mkDebugOperation(mod_3047_inner, "mod_3047");
    Operation_IFC mod_3048_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3048 <- mkDebugOperation(mod_3048_inner, "mod_3048");
    Operation_IFC mod_3049_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3049 <- mkDebugOperation(mod_3049_inner, "mod_3049");
    Operation_IFC mod_3050_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3050 <- mkDebugOperation(mod_3050_inner, "mod_3050");
    Operation_IFC mod_3051_inner <- mkBinaryMap(2749, mul_tile);
    Operation_IFC mod_3051 <- mkDebugOperation(mod_3051_inner, "mod_3051");
    PMU_IFC mod_3052_bufferize <- mkPMU(1);
    Operation_IFC mod_3052_inner = mod_3052_bufferize.operation;
    Operation_IFC mod_3052 <- mkDebugOperation(mod_3052_inner, "mod_3052");
    PMU_IFC mod_3053_bufferize <- mkPMU(2);
    Operation_IFC mod_3053_inner = mod_3053_bufferize.operation;
    Operation_IFC mod_3053 <- mkDebugOperation(mod_3053_inner, "mod_3053");
    PMU_IFC mod_3054_bufferize <- mkPMU(2);
    Operation_IFC mod_3054_inner = mod_3054_bufferize.operation;
    Operation_IFC mod_3054 <- mkDebugOperation(mod_3054_inner, "mod_3054");
    Operation_IFC mod_3055_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3055 <- mkDebugOperation(mod_3055_inner, "mod_3055");
    Operation_IFC mod_3056_inner <- mkFlatten(1);
    Operation_IFC mod_3056 <- mkDebugOperation(mod_3056_inner, "mod_3056");
    Operation_IFC mod_3057_inner <- mkFlatten(0);
    Operation_IFC mod_3057 <- mkDebugOperation(mod_3057_inner, "mod_3057");
    Operation_IFC mod_3058_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3058 <- mkDebugOperation(mod_3058_inner, "mod_3058");
    Operation_IFC mod_3059_inner <- mkUnaryMap(1722, silu_tile);
    Operation_IFC mod_3059 <- mkDebugOperation(mod_3059_inner, "mod_3059");
    Operation_IFC mod_3060_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3060 <- mkDebugOperation(mod_3060_inner, "mod_3060");
    Operation_IFC mod_3061_inner <- mkBinaryMap(1594, matmul_t_tile);
    Operation_IFC mod_3061 <- mkDebugOperation(mod_3061_inner, "mod_3061");
    PMU_IFC mod_3062_bufferize <- mkPMU(2);
    Operation_IFC mod_3062_inner = mod_3062_bufferize.operation;
    Operation_IFC mod_3062 <- mkDebugOperation(mod_3062_inner, "mod_3062");
    Operation_IFC mod_3063_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3063 <- mkDebugOperation(mod_3063_inner, "mod_3063");
    Operation_IFC mod_3064_inner <- mkFlatten(1);
    Operation_IFC mod_3064 <- mkDebugOperation(mod_3064_inner, "mod_3064");
    Operation_IFC mod_3065_inner <- mkFlatten(0);
    Operation_IFC mod_3065 <- mkDebugOperation(mod_3065_inner, "mod_3065");
    PMU_IFC mod_3066_bufferize <- mkPMU(1);
    Operation_IFC mod_3066_inner = mod_3066_bufferize.operation;
    Operation_IFC mod_3066 <- mkDebugOperation(mod_3066_inner, "mod_3066");
    Operation_IFC mod_3067_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3067 <- mkDebugOperation(mod_3067_inner, "mod_3067");
    PMU_IFC mod_3068_bufferize <- mkPMU(2);
    Operation_IFC mod_3068_inner = mod_3068_bufferize.operation;
    Operation_IFC mod_3068 <- mkDebugOperation(mod_3068_inner, "mod_3068");
    Operation_IFC mod_3069_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3069 <- mkDebugOperation(mod_3069_inner, "mod_3069");
    Operation_IFC mod_3070_inner <- mkFlatten(1);
    Operation_IFC mod_3070 <- mkDebugOperation(mod_3070_inner, "mod_3070");
    Operation_IFC mod_3071_inner <- mkFlatten(0);
    Operation_IFC mod_3071 <- mkDebugOperation(mod_3071_inner, "mod_3071");
    Operation_IFC mod_3072_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3072 <- mkDebugOperation(mod_3072_inner, "mod_3072");
    Operation_IFC mod_3073_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3073 <- mkDebugOperation(mod_3073_inner, "mod_3073");
    PMU_IFC mod_3074_bufferize <- mkPMU(2);
    Operation_IFC mod_3074_inner = mod_3074_bufferize.operation;
    Operation_IFC mod_3074 <- mkDebugOperation(mod_3074_inner, "mod_3074");
    rule rule_3923;
        ChannelMessage t;
        t <- mod_3035.get(0);
        mod_3036.put(0, t);
    endrule
    rule rule_3924;
        ChannelMessage t;
        t <- mod_3061.get(0);
        mod_3060.put(0, t);
    endrule
    rule rule_3925;
        ChannelMessage t;
        t <- mod_3060.get(0);
        mod_3059.put(0, t);
    endrule
    rule rule_3926;
        ChannelMessage t;
        t <- mod_3066.get(0);
        mod_3067.put(0, t);
    endrule
    rule rule_3927;
        ChannelMessage t;
        t <- mod_3058.get(0);
        mod_3046.put(1, t);
    endrule
    rule rule_3928;
        ChannelMessage t;
        t <- mod_3062.get(0);
        mod_3063.put(0, t);
    endrule
    rule rule_3929;
        ChannelMessage t;
        t <- mod_3069.get(0);
        mod_3068.put(1, t);
    endrule
    rule rule_3930;
        ChannelMessage t;
        t <- mod_3042.get(0);
        mod_3072.put(0, t);
    endrule
    rule rule_3931;
        ChannelMessage t;
        t <- mod_3041.get(1);
        mod_3042.put(0, t);
    endrule
    rule rule_3932;
        ChannelMessage t;
        t <- mod_3050.get(0);
        mod_3052.put(0, t);
    endrule
    rule rule_3933;
        ChannelMessage t;
        t <- mod_3053.get(0);
        mod_3053.put(1, t);
    endrule
    rule rule_3934;
        ChannelMessage t;
        t <- mod_3063.get(0);
        mod_3062.put(1, t);
    endrule
    rule rule_3935;
        ChannelMessage t;
        t <- mod_3046.get(0);
        mod_3058.put(0, t);
    endrule
    rule rule_3936;
        ChannelMessage t;
        t <- mod_3052.get(1);
        mod_3050.put(1, t);
    endrule
    rule rule_3937;
        ChannelMessage t;
        t <- mod_3067.get(0);
        mod_3066.put(1, t);
    endrule
    rule rule_3938;
        ChannelMessage t;
        t <- mod_3071.get(0);
        mod_3070.put(0, t);
    endrule
    rule rule_3939;
        ChannelMessage t;
        t <- mod_3053.get(1);
        mod_3049.put(1, t);
    endrule
    rule rule_3940;
        ChannelMessage t;
        t <- mod_3056.get(0);
        mod_3054.put(0, t);
    endrule
    rule rule_3941;
        ChannelMessage t;
        t <- mod_3062.get(1);
        mod_3061.put(1, t);
    endrule
    rule rule_3942;
        ChannelMessage t;
        t <- mod_3043.get(0);
        mod_3044.put(0, t);
    endrule
    rule rule_3943;
        ChannelMessage t;
        t <- mod_3042.get(1);
        mod_3043.put(0, t);
    endrule
    rule rule_3944;
        ChannelMessage t;
        t <- mod_3039.get(3);
        mod_3040.put(0, t);
    endrule
    rule rule_3945;
        ChannelMessage t;
        t <- mod_3074.get(1);
        mod_3038.put(1, t);
    endrule
    rule rule_3946;
        ChannelMessage t;
        t <- mod_3054.get(0);
        mod_3055.put(0, t);
    endrule
    rule rule_3947;
        ChannelMessage t;
        t <- mod_3074.get(0);
        mod_3074.put(1, t);
    endrule
    rule rule_3948;
        ChannelMessage t;
        t <- mod_3046.get(1);
        mod_3047.put(0, t);
    endrule
    rule rule_3949;
        ChannelMessage t;
        t <- mod_3038.get(1);
        mod_3039.put(0, t);
    endrule
    rule rule_3950;
        ChannelMessage t;
        t <- mod_3045.get(0);
        mod_3046.put(0, t);
    endrule
    rule rule_3951;
        ChannelMessage t;
        t <- mod_3037.get(0);
        mod_3038.put(0, t);
    endrule
    rule rule_3952;
        ChannelMessage t;
        t <- mod_3057.get(0);
        mod_3056.put(0, t);
    endrule
    rule rule_3953;
        ChannelMessage t;
        t <- mod_3049.get(0);
        mod_3053.put(0, t);
    endrule
    rule rule_3954;
        ChannelMessage t;
        t <- mod_3040.get(1);
        mod_3041.put(0, t);
    endrule
    rule rule_3955;
        ChannelMessage t;
        t <- mod_3052.get(0);
        mod_3052.put(1, t);
    endrule
    rule rule_3956;
        ChannelMessage t;
        t <- mod_3036.get(0);
        mod_3037.put(0, t);
    endrule
    rule rule_3957;
        ChannelMessage t;
        t <- mod_3064.get(0);
        mod_3062.put(0, t);
    endrule
    rule rule_3958;
        ChannelMessage t;
        t <- mod_3072.get(0);
        mod_3042.put(1, t);
    endrule
    rule rule_3959;
        ChannelMessage t;
        t <- mod_3038.get(0);
        mod_3074.put(0, t);
    endrule
    rule rule_3960;
        ChannelMessage t;
        t <- mod_3049.get(1);
        mod_3050.put(0, t);
    endrule
    rule rule_3961;
        ChannelMessage t;
        t <- mod_3044.get(0);
        mod_3045.put(0, t);
    endrule
    rule rule_3962;
        ChannelMessage t;
        t <- mod_3066.get(1);
        mod_3061.put(0, t);
    endrule
    rule rule_3963;
        ChannelMessage t;
        t <- mod_3065.get(0);
        mod_3064.put(0, t);
    endrule
    rule rule_3964;
        ChannelMessage t;
        t <- mod_3041.get(0);
        mod_3066.put(0, t);
    endrule
    rule rule_3965;
        ChannelMessage t;
        t <- mod_3059.get(0);
        mod_3045.put(1, t);
    endrule
    rule rule_3966;
        ChannelMessage t;
        t <- mod_3070.get(0);
        mod_3068.put(0, t);
    endrule
    rule rule_3967;
        ChannelMessage t;
        t <- mod_3054.get(1);
        mod_3047.put(1, t);
    endrule
    rule rule_3968;
        ChannelMessage t;
        t <- mod_3055.get(0);
        mod_3054.put(1, t);
    endrule
    rule rule_3969;
        ChannelMessage t;
        t <- mod_3068.get(0);
        mod_3069.put(0, t);
    endrule
    rule rule_3970;
        ChannelMessage t;
        t <- mod_3040.get(0);
        mod_3073.put(0, t);
    endrule
    rule rule_3971;
        ChannelMessage t;
        t <- mod_3050.get(1);
        mod_3051.put(1, t);
    endrule
    rule rule_3972;
        ChannelMessage t;
        t <- mod_3068.get(1);
        mod_3043.put(1, t);
    endrule
    rule rule_3973;
        ChannelMessage t;
        t <- mod_3073.get(0);
        mod_3040.put(1, t);
    endrule
    rule rule_3974;
        ChannelMessage t;
        t <- mod_3047.get(0);
        mod_3048.put(0, t);
    endrule
    rule rule_3975;
        ChannelMessage t;
        t <- mod_3048.get(0);
        mod_3049.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3035.put(0, t);
        end
        if (i == 1) begin
            mod_3051.put(0, t);
        end
        if (i == 2) begin
            mod_3057.put(0, t);
        end
        if (i == 3) begin
            mod_3065.put(0, t);
        end
        if (i == 4) begin
            mod_3071.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 2) begin
            t <- mod_3039.get(0);
        end
        if (i == 1) begin
            t <- mod_3039.get(1);
        end
        if (i == 3) begin
            t <- mod_3039.get(2);
        end
        if (i == 0) begin
            t <- mod_3051.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6109 (Operation_IFC);
    Operation_IFC mod_3076_inner <- mkReshape(2, 64);
    Operation_IFC mod_3076 <- mkDebugOperation(mod_3076_inner, "mod_3076");
    Operation_IFC mod_3077_inner <- mkFlatten(1);
    Operation_IFC mod_3077 <- mkDebugOperation(mod_3077_inner, "mod_3077");
    Operation_IFC mod_3078_inner <- mkFlatten(2);
    Operation_IFC mod_3078 <- mkDebugOperation(mod_3078_inner, "mod_3078");
    Operation_IFC mod_3079_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3079 <- mkDebugOperation(mod_3079_inner, "mod_3079");
    Broadcast_IFC#(4) mod_3080_inner <- mkBroadcast(4);
    Operation_IFC mod_3080 <- mkDebugOperation(mod_3080_inner.op, "mod_3080");
    PMU_IFC mod_3081_bufferize <- mkPMU(2);
    Operation_IFC mod_3081_inner = mod_3081_bufferize.operation;
    Operation_IFC mod_3081 <- mkDebugOperation(mod_3081_inner, "mod_3081");
    Broadcast_IFC#(2) mod_3082_inner <- mkBroadcast(2);
    Operation_IFC mod_3082 <- mkDebugOperation(mod_3082_inner.op, "mod_3082");
    PMU_IFC mod_3083_bufferize <- mkPMU(1);
    Operation_IFC mod_3083_inner = mod_3083_bufferize.operation;
    Operation_IFC mod_3083 <- mkDebugOperation(mod_3083_inner, "mod_3083");
    Operation_IFC mod_3084_inner <- mkBinaryMap(1081, matmul_t_tile);
    Operation_IFC mod_3084 <- mkDebugOperation(mod_3084_inner, "mod_3084");
    Operation_IFC mod_3085_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3085 <- mkDebugOperation(mod_3085_inner, "mod_3085");
    Operation_IFC mod_3086_inner <- mkBinaryMap(1849, mul_tile);
    Operation_IFC mod_3086 <- mkDebugOperation(mod_3086_inner, "mod_3086");
    PMU_IFC mod_3087_bufferize <- mkPMU(1);
    Operation_IFC mod_3087_inner = mod_3087_bufferize.operation;
    Operation_IFC mod_3087 <- mkDebugOperation(mod_3087_inner, "mod_3087");
    Operation_IFC mod_3088_inner <- mkBinaryMap(2413, matmul_t_tile);
    Operation_IFC mod_3088 <- mkDebugOperation(mod_3088_inner, "mod_3088");
    Operation_IFC mod_3089_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3089 <- mkDebugOperation(mod_3089_inner, "mod_3089");
    Operation_IFC mod_3090_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3090 <- mkDebugOperation(mod_3090_inner, "mod_3090");
    Operation_IFC mod_3091_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3091 <- mkDebugOperation(mod_3091_inner, "mod_3091");
    Operation_IFC mod_3092_inner <- mkBinaryMap(2748, mul_tile);
    Operation_IFC mod_3092 <- mkDebugOperation(mod_3092_inner, "mod_3092");
    PMU_IFC mod_3093_bufferize <- mkPMU(1);
    Operation_IFC mod_3093_inner = mod_3093_bufferize.operation;
    Operation_IFC mod_3093 <- mkDebugOperation(mod_3093_inner, "mod_3093");
    PMU_IFC mod_3094_bufferize <- mkPMU(2);
    Operation_IFC mod_3094_inner = mod_3094_bufferize.operation;
    Operation_IFC mod_3094 <- mkDebugOperation(mod_3094_inner, "mod_3094");
    PMU_IFC mod_3095_bufferize <- mkPMU(2);
    Operation_IFC mod_3095_inner = mod_3095_bufferize.operation;
    Operation_IFC mod_3095 <- mkDebugOperation(mod_3095_inner, "mod_3095");
    Operation_IFC mod_3096_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3096 <- mkDebugOperation(mod_3096_inner, "mod_3096");
    Operation_IFC mod_3097_inner <- mkFlatten(1);
    Operation_IFC mod_3097 <- mkDebugOperation(mod_3097_inner, "mod_3097");
    Operation_IFC mod_3098_inner <- mkFlatten(0);
    Operation_IFC mod_3098 <- mkDebugOperation(mod_3098_inner, "mod_3098");
    Operation_IFC mod_3099_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3099 <- mkDebugOperation(mod_3099_inner, "mod_3099");
    Operation_IFC mod_3100_inner <- mkUnaryMap(1721, silu_tile);
    Operation_IFC mod_3100 <- mkDebugOperation(mod_3100_inner, "mod_3100");
    Operation_IFC mod_3101_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3101 <- mkDebugOperation(mod_3101_inner, "mod_3101");
    Operation_IFC mod_3102_inner <- mkBinaryMap(1593, matmul_t_tile);
    Operation_IFC mod_3102 <- mkDebugOperation(mod_3102_inner, "mod_3102");
    PMU_IFC mod_3103_bufferize <- mkPMU(2);
    Operation_IFC mod_3103_inner = mod_3103_bufferize.operation;
    Operation_IFC mod_3103 <- mkDebugOperation(mod_3103_inner, "mod_3103");
    Operation_IFC mod_3104_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3104 <- mkDebugOperation(mod_3104_inner, "mod_3104");
    Operation_IFC mod_3105_inner <- mkFlatten(1);
    Operation_IFC mod_3105 <- mkDebugOperation(mod_3105_inner, "mod_3105");
    Operation_IFC mod_3106_inner <- mkFlatten(0);
    Operation_IFC mod_3106 <- mkDebugOperation(mod_3106_inner, "mod_3106");
    PMU_IFC mod_3107_bufferize <- mkPMU(1);
    Operation_IFC mod_3107_inner = mod_3107_bufferize.operation;
    Operation_IFC mod_3107 <- mkDebugOperation(mod_3107_inner, "mod_3107");
    Operation_IFC mod_3108_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3108 <- mkDebugOperation(mod_3108_inner, "mod_3108");
    PMU_IFC mod_3109_bufferize <- mkPMU(2);
    Operation_IFC mod_3109_inner = mod_3109_bufferize.operation;
    Operation_IFC mod_3109 <- mkDebugOperation(mod_3109_inner, "mod_3109");
    Operation_IFC mod_3110_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3110 <- mkDebugOperation(mod_3110_inner, "mod_3110");
    Operation_IFC mod_3111_inner <- mkFlatten(1);
    Operation_IFC mod_3111 <- mkDebugOperation(mod_3111_inner, "mod_3111");
    Operation_IFC mod_3112_inner <- mkFlatten(0);
    Operation_IFC mod_3112 <- mkDebugOperation(mod_3112_inner, "mod_3112");
    Operation_IFC mod_3113_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3113 <- mkDebugOperation(mod_3113_inner, "mod_3113");
    Operation_IFC mod_3114_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3114 <- mkDebugOperation(mod_3114_inner, "mod_3114");
    PMU_IFC mod_3115_bufferize <- mkPMU(2);
    Operation_IFC mod_3115_inner = mod_3115_bufferize.operation;
    Operation_IFC mod_3115 <- mkDebugOperation(mod_3115_inner, "mod_3115");
    rule rule_3976;
        ChannelMessage t;
        t <- mod_3084.get(0);
        mod_3085.put(0, t);
    endrule
    rule rule_3977;
        ChannelMessage t;
        t <- mod_3108.get(0);
        mod_3107.put(1, t);
    endrule
    rule rule_3978;
        ChannelMessage t;
        t <- mod_3079.get(0);
        mod_3115.put(0, t);
    endrule
    rule rule_3979;
        ChannelMessage t;
        t <- mod_3094.get(0);
        mod_3094.put(1, t);
    endrule
    rule rule_3980;
        ChannelMessage t;
        t <- mod_3078.get(0);
        mod_3079.put(0, t);
    endrule
    rule rule_3981;
        ChannelMessage t;
        t <- mod_3079.get(1);
        mod_3080.put(0, t);
    endrule
    rule rule_3982;
        ChannelMessage t;
        t <- mod_3103.get(1);
        mod_3102.put(1, t);
    endrule
    rule rule_3983;
        ChannelMessage t;
        t <- mod_3100.get(0);
        mod_3086.put(1, t);
    endrule
    rule rule_3984;
        ChannelMessage t;
        t <- mod_3106.get(0);
        mod_3105.put(0, t);
    endrule
    rule rule_3985;
        ChannelMessage t;
        t <- mod_3096.get(0);
        mod_3095.put(1, t);
    endrule
    rule rule_3986;
        ChannelMessage t;
        t <- mod_3115.get(0);
        mod_3115.put(1, t);
    endrule
    rule rule_3987;
        ChannelMessage t;
        t <- mod_3090.get(0);
        mod_3094.put(0, t);
    endrule
    rule rule_3988;
        ChannelMessage t;
        t <- mod_3094.get(1);
        mod_3090.put(1, t);
    endrule
    rule rule_3989;
        ChannelMessage t;
        t <- mod_3091.get(0);
        mod_3093.put(0, t);
    endrule
    rule rule_3990;
        ChannelMessage t;
        t <- mod_3087.get(0);
        mod_3099.put(0, t);
    endrule
    rule rule_3991;
        ChannelMessage t;
        t <- mod_3088.get(0);
        mod_3089.put(0, t);
    endrule
    rule rule_3992;
        ChannelMessage t;
        t <- mod_3093.get(0);
        mod_3093.put(1, t);
    endrule
    rule rule_3993;
        ChannelMessage t;
        t <- mod_3107.get(1);
        mod_3102.put(0, t);
    endrule
    rule rule_3994;
        ChannelMessage t;
        t <- mod_3115.get(1);
        mod_3079.put(1, t);
    endrule
    rule rule_3995;
        ChannelMessage t;
        t <- mod_3090.get(1);
        mod_3091.put(0, t);
    endrule
    rule rule_3996;
        ChannelMessage t;
        t <- mod_3086.get(0);
        mod_3087.put(0, t);
    endrule
    rule rule_3997;
        ChannelMessage t;
        t <- mod_3087.get(1);
        mod_3088.put(0, t);
    endrule
    rule rule_3998;
        ChannelMessage t;
        t <- mod_3083.get(0);
        mod_3113.put(0, t);
    endrule
    rule rule_3999;
        ChannelMessage t;
        t <- mod_3109.get(1);
        mod_3084.put(1, t);
    endrule
    rule rule_4000;
        ChannelMessage t;
        t <- mod_3077.get(0);
        mod_3078.put(0, t);
    endrule
    rule rule_4001;
        ChannelMessage t;
        t <- mod_3103.get(0);
        mod_3104.put(0, t);
    endrule
    rule rule_4002;
        ChannelMessage t;
        t <- mod_3101.get(0);
        mod_3100.put(0, t);
    endrule
    rule rule_4003;
        ChannelMessage t;
        t <- mod_3089.get(0);
        mod_3090.put(0, t);
    endrule
    rule rule_4004;
        ChannelMessage t;
        t <- mod_3082.get(0);
        mod_3107.put(0, t);
    endrule
    rule rule_4005;
        ChannelMessage t;
        t <- mod_3085.get(0);
        mod_3086.put(0, t);
    endrule
    rule rule_4006;
        ChannelMessage t;
        t <- mod_3080.get(3);
        mod_3081.put(0, t);
    endrule
    rule rule_4007;
        ChannelMessage t;
        t <- mod_3083.get(1);
        mod_3084.put(0, t);
    endrule
    rule rule_4008;
        ChannelMessage t;
        t <- mod_3109.get(0);
        mod_3110.put(0, t);
    endrule
    rule rule_4009;
        ChannelMessage t;
        t <- mod_3105.get(0);
        mod_3103.put(0, t);
    endrule
    rule rule_4010;
        ChannelMessage t;
        t <- mod_3081.get(1);
        mod_3082.put(0, t);
    endrule
    rule rule_4011;
        ChannelMessage t;
        t <- mod_3104.get(0);
        mod_3103.put(1, t);
    endrule
    rule rule_4012;
        ChannelMessage t;
        t <- mod_3113.get(0);
        mod_3083.put(1, t);
    endrule
    rule rule_4013;
        ChannelMessage t;
        t <- mod_3114.get(0);
        mod_3081.put(1, t);
    endrule
    rule rule_4014;
        ChannelMessage t;
        t <- mod_3081.get(0);
        mod_3114.put(0, t);
    endrule
    rule rule_4015;
        ChannelMessage t;
        t <- mod_3082.get(1);
        mod_3083.put(0, t);
    endrule
    rule rule_4016;
        ChannelMessage t;
        t <- mod_3091.get(1);
        mod_3092.put(1, t);
    endrule
    rule rule_4017;
        ChannelMessage t;
        t <- mod_3107.get(0);
        mod_3108.put(0, t);
    endrule
    rule rule_4018;
        ChannelMessage t;
        t <- mod_3095.get(1);
        mod_3088.put(1, t);
    endrule
    rule rule_4019;
        ChannelMessage t;
        t <- mod_3093.get(1);
        mod_3091.put(1, t);
    endrule
    rule rule_4020;
        ChannelMessage t;
        t <- mod_3095.get(0);
        mod_3096.put(0, t);
    endrule
    rule rule_4021;
        ChannelMessage t;
        t <- mod_3097.get(0);
        mod_3095.put(0, t);
    endrule
    rule rule_4022;
        ChannelMessage t;
        t <- mod_3112.get(0);
        mod_3111.put(0, t);
    endrule
    rule rule_4023;
        ChannelMessage t;
        t <- mod_3098.get(0);
        mod_3097.put(0, t);
    endrule
    rule rule_4024;
        ChannelMessage t;
        t <- mod_3076.get(0);
        mod_3077.put(0, t);
    endrule
    rule rule_4025;
        ChannelMessage t;
        t <- mod_3099.get(0);
        mod_3087.put(1, t);
    endrule
    rule rule_4026;
        ChannelMessage t;
        t <- mod_3110.get(0);
        mod_3109.put(1, t);
    endrule
    rule rule_4027;
        ChannelMessage t;
        t <- mod_3111.get(0);
        mod_3109.put(0, t);
    endrule
    rule rule_4028;
        ChannelMessage t;
        t <- mod_3102.get(0);
        mod_3101.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3076.put(0, t);
        end
        if (i == 1) begin
            mod_3092.put(0, t);
        end
        if (i == 2) begin
            mod_3098.put(0, t);
        end
        if (i == 3) begin
            mod_3106.put(0, t);
        end
        if (i == 4) begin
            mod_3112.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_3080.get(0);
        end
        if (i == 2) begin
            t <- mod_3080.get(1);
        end
        if (i == 0) begin
            t <- mod_3080.get(2);
        end
        if (i == 1) begin
            t <- mod_3092.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6110 (Operation_IFC);
    Operation_IFC mod_3117_inner <- mkReshape(2, 64);
    Operation_IFC mod_3117 <- mkDebugOperation(mod_3117_inner, "mod_3117");
    Operation_IFC mod_3118_inner <- mkFlatten(1);
    Operation_IFC mod_3118 <- mkDebugOperation(mod_3118_inner, "mod_3118");
    Operation_IFC mod_3119_inner <- mkFlatten(2);
    Operation_IFC mod_3119 <- mkDebugOperation(mod_3119_inner, "mod_3119");
    Operation_IFC mod_3120_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3120 <- mkDebugOperation(mod_3120_inner, "mod_3120");
    Broadcast_IFC#(4) mod_3121_inner <- mkBroadcast(4);
    Operation_IFC mod_3121 <- mkDebugOperation(mod_3121_inner.op, "mod_3121");
    PMU_IFC mod_3122_bufferize <- mkPMU(2);
    Operation_IFC mod_3122_inner = mod_3122_bufferize.operation;
    Operation_IFC mod_3122 <- mkDebugOperation(mod_3122_inner, "mod_3122");
    Broadcast_IFC#(2) mod_3123_inner <- mkBroadcast(2);
    Operation_IFC mod_3123 <- mkDebugOperation(mod_3123_inner.op, "mod_3123");
    PMU_IFC mod_3124_bufferize <- mkPMU(1);
    Operation_IFC mod_3124_inner = mod_3124_bufferize.operation;
    Operation_IFC mod_3124 <- mkDebugOperation(mod_3124_inner, "mod_3124");
    Operation_IFC mod_3125_inner <- mkBinaryMap(1080, matmul_t_tile);
    Operation_IFC mod_3125 <- mkDebugOperation(mod_3125_inner, "mod_3125");
    Operation_IFC mod_3126_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3126 <- mkDebugOperation(mod_3126_inner, "mod_3126");
    Operation_IFC mod_3127_inner <- mkBinaryMap(1848, mul_tile);
    Operation_IFC mod_3127 <- mkDebugOperation(mod_3127_inner, "mod_3127");
    PMU_IFC mod_3128_bufferize <- mkPMU(1);
    Operation_IFC mod_3128_inner = mod_3128_bufferize.operation;
    Operation_IFC mod_3128 <- mkDebugOperation(mod_3128_inner, "mod_3128");
    Operation_IFC mod_3129_inner <- mkBinaryMap(2411, matmul_t_tile);
    Operation_IFC mod_3129 <- mkDebugOperation(mod_3129_inner, "mod_3129");
    Operation_IFC mod_3130_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3130 <- mkDebugOperation(mod_3130_inner, "mod_3130");
    Operation_IFC mod_3131_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3131 <- mkDebugOperation(mod_3131_inner, "mod_3131");
    Operation_IFC mod_3132_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3132 <- mkDebugOperation(mod_3132_inner, "mod_3132");
    Operation_IFC mod_3133_inner <- mkBinaryMap(2747, mul_tile);
    Operation_IFC mod_3133 <- mkDebugOperation(mod_3133_inner, "mod_3133");
    PMU_IFC mod_3134_bufferize <- mkPMU(1);
    Operation_IFC mod_3134_inner = mod_3134_bufferize.operation;
    Operation_IFC mod_3134 <- mkDebugOperation(mod_3134_inner, "mod_3134");
    PMU_IFC mod_3135_bufferize <- mkPMU(2);
    Operation_IFC mod_3135_inner = mod_3135_bufferize.operation;
    Operation_IFC mod_3135 <- mkDebugOperation(mod_3135_inner, "mod_3135");
    PMU_IFC mod_3136_bufferize <- mkPMU(2);
    Operation_IFC mod_3136_inner = mod_3136_bufferize.operation;
    Operation_IFC mod_3136 <- mkDebugOperation(mod_3136_inner, "mod_3136");
    Operation_IFC mod_3137_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3137 <- mkDebugOperation(mod_3137_inner, "mod_3137");
    Operation_IFC mod_3138_inner <- mkFlatten(1);
    Operation_IFC mod_3138 <- mkDebugOperation(mod_3138_inner, "mod_3138");
    Operation_IFC mod_3139_inner <- mkFlatten(0);
    Operation_IFC mod_3139 <- mkDebugOperation(mod_3139_inner, "mod_3139");
    Operation_IFC mod_3140_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3140 <- mkDebugOperation(mod_3140_inner, "mod_3140");
    Operation_IFC mod_3141_inner <- mkUnaryMap(1720, silu_tile);
    Operation_IFC mod_3141 <- mkDebugOperation(mod_3141_inner, "mod_3141");
    Operation_IFC mod_3142_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3142 <- mkDebugOperation(mod_3142_inner, "mod_3142");
    Operation_IFC mod_3143_inner <- mkBinaryMap(1592, matmul_t_tile);
    Operation_IFC mod_3143 <- mkDebugOperation(mod_3143_inner, "mod_3143");
    PMU_IFC mod_3144_bufferize <- mkPMU(2);
    Operation_IFC mod_3144_inner = mod_3144_bufferize.operation;
    Operation_IFC mod_3144 <- mkDebugOperation(mod_3144_inner, "mod_3144");
    Operation_IFC mod_3145_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3145 <- mkDebugOperation(mod_3145_inner, "mod_3145");
    Operation_IFC mod_3146_inner <- mkFlatten(1);
    Operation_IFC mod_3146 <- mkDebugOperation(mod_3146_inner, "mod_3146");
    Operation_IFC mod_3147_inner <- mkFlatten(0);
    Operation_IFC mod_3147 <- mkDebugOperation(mod_3147_inner, "mod_3147");
    PMU_IFC mod_3148_bufferize <- mkPMU(1);
    Operation_IFC mod_3148_inner = mod_3148_bufferize.operation;
    Operation_IFC mod_3148 <- mkDebugOperation(mod_3148_inner, "mod_3148");
    Operation_IFC mod_3149_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3149 <- mkDebugOperation(mod_3149_inner, "mod_3149");
    PMU_IFC mod_3150_bufferize <- mkPMU(2);
    Operation_IFC mod_3150_inner = mod_3150_bufferize.operation;
    Operation_IFC mod_3150 <- mkDebugOperation(mod_3150_inner, "mod_3150");
    Operation_IFC mod_3151_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3151 <- mkDebugOperation(mod_3151_inner, "mod_3151");
    Operation_IFC mod_3152_inner <- mkFlatten(1);
    Operation_IFC mod_3152 <- mkDebugOperation(mod_3152_inner, "mod_3152");
    Operation_IFC mod_3153_inner <- mkFlatten(0);
    Operation_IFC mod_3153 <- mkDebugOperation(mod_3153_inner, "mod_3153");
    Operation_IFC mod_3154_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3154 <- mkDebugOperation(mod_3154_inner, "mod_3154");
    Operation_IFC mod_3155_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3155 <- mkDebugOperation(mod_3155_inner, "mod_3155");
    PMU_IFC mod_3156_bufferize <- mkPMU(2);
    Operation_IFC mod_3156_inner = mod_3156_bufferize.operation;
    Operation_IFC mod_3156 <- mkDebugOperation(mod_3156_inner, "mod_3156");
    rule rule_4029;
        ChannelMessage t;
        t <- mod_3150.get(1);
        mod_3125.put(1, t);
    endrule
    rule rule_4030;
        ChannelMessage t;
        t <- mod_3128.get(0);
        mod_3140.put(0, t);
    endrule
    rule rule_4031;
        ChannelMessage t;
        t <- mod_3128.get(1);
        mod_3129.put(0, t);
    endrule
    rule rule_4032;
        ChannelMessage t;
        t <- mod_3123.get(0);
        mod_3148.put(0, t);
    endrule
    rule rule_4033;
        ChannelMessage t;
        t <- mod_3152.get(0);
        mod_3150.put(0, t);
    endrule
    rule rule_4034;
        ChannelMessage t;
        t <- mod_3155.get(0);
        mod_3122.put(1, t);
    endrule
    rule rule_4035;
        ChannelMessage t;
        t <- mod_3132.get(1);
        mod_3133.put(1, t);
    endrule
    rule rule_4036;
        ChannelMessage t;
        t <- mod_3149.get(0);
        mod_3148.put(1, t);
    endrule
    rule rule_4037;
        ChannelMessage t;
        t <- mod_3153.get(0);
        mod_3152.put(0, t);
    endrule
    rule rule_4038;
        ChannelMessage t;
        t <- mod_3125.get(0);
        mod_3126.put(0, t);
    endrule
    rule rule_4039;
        ChannelMessage t;
        t <- mod_3135.get(1);
        mod_3131.put(1, t);
    endrule
    rule rule_4040;
        ChannelMessage t;
        t <- mod_3123.get(1);
        mod_3124.put(0, t);
    endrule
    rule rule_4041;
        ChannelMessage t;
        t <- mod_3154.get(0);
        mod_3124.put(1, t);
    endrule
    rule rule_4042;
        ChannelMessage t;
        t <- mod_3124.get(1);
        mod_3125.put(0, t);
    endrule
    rule rule_4043;
        ChannelMessage t;
        t <- mod_3121.get(3);
        mod_3122.put(0, t);
    endrule
    rule rule_4044;
        ChannelMessage t;
        t <- mod_3118.get(0);
        mod_3119.put(0, t);
    endrule
    rule rule_4045;
        ChannelMessage t;
        t <- mod_3150.get(0);
        mod_3151.put(0, t);
    endrule
    rule rule_4046;
        ChannelMessage t;
        t <- mod_3136.get(0);
        mod_3137.put(0, t);
    endrule
    rule rule_4047;
        ChannelMessage t;
        t <- mod_3144.get(0);
        mod_3145.put(0, t);
    endrule
    rule rule_4048;
        ChannelMessage t;
        t <- mod_3129.get(0);
        mod_3130.put(0, t);
    endrule
    rule rule_4049;
        ChannelMessage t;
        t <- mod_3122.get(0);
        mod_3155.put(0, t);
    endrule
    rule rule_4050;
        ChannelMessage t;
        t <- mod_3120.get(0);
        mod_3156.put(0, t);
    endrule
    rule rule_4051;
        ChannelMessage t;
        t <- mod_3131.get(1);
        mod_3132.put(0, t);
    endrule
    rule rule_4052;
        ChannelMessage t;
        t <- mod_3137.get(0);
        mod_3136.put(1, t);
    endrule
    rule rule_4053;
        ChannelMessage t;
        t <- mod_3132.get(0);
        mod_3134.put(0, t);
    endrule
    rule rule_4054;
        ChannelMessage t;
        t <- mod_3130.get(0);
        mod_3131.put(0, t);
    endrule
    rule rule_4055;
        ChannelMessage t;
        t <- mod_3142.get(0);
        mod_3141.put(0, t);
    endrule
    rule rule_4056;
        ChannelMessage t;
        t <- mod_3126.get(0);
        mod_3127.put(0, t);
    endrule
    rule rule_4057;
        ChannelMessage t;
        t <- mod_3145.get(0);
        mod_3144.put(1, t);
    endrule
    rule rule_4058;
        ChannelMessage t;
        t <- mod_3124.get(0);
        mod_3154.put(0, t);
    endrule
    rule rule_4059;
        ChannelMessage t;
        t <- mod_3117.get(0);
        mod_3118.put(0, t);
    endrule
    rule rule_4060;
        ChannelMessage t;
        t <- mod_3119.get(0);
        mod_3120.put(0, t);
    endrule
    rule rule_4061;
        ChannelMessage t;
        t <- mod_3134.get(0);
        mod_3134.put(1, t);
    endrule
    rule rule_4062;
        ChannelMessage t;
        t <- mod_3141.get(0);
        mod_3127.put(1, t);
    endrule
    rule rule_4063;
        ChannelMessage t;
        t <- mod_3122.get(1);
        mod_3123.put(0, t);
    endrule
    rule rule_4064;
        ChannelMessage t;
        t <- mod_3144.get(1);
        mod_3143.put(1, t);
    endrule
    rule rule_4065;
        ChannelMessage t;
        t <- mod_3131.get(0);
        mod_3135.put(0, t);
    endrule
    rule rule_4066;
        ChannelMessage t;
        t <- mod_3146.get(0);
        mod_3144.put(0, t);
    endrule
    rule rule_4067;
        ChannelMessage t;
        t <- mod_3147.get(0);
        mod_3146.put(0, t);
    endrule
    rule rule_4068;
        ChannelMessage t;
        t <- mod_3136.get(1);
        mod_3129.put(1, t);
    endrule
    rule rule_4069;
        ChannelMessage t;
        t <- mod_3140.get(0);
        mod_3128.put(1, t);
    endrule
    rule rule_4070;
        ChannelMessage t;
        t <- mod_3138.get(0);
        mod_3136.put(0, t);
    endrule
    rule rule_4071;
        ChannelMessage t;
        t <- mod_3139.get(0);
        mod_3138.put(0, t);
    endrule
    rule rule_4072;
        ChannelMessage t;
        t <- mod_3143.get(0);
        mod_3142.put(0, t);
    endrule
    rule rule_4073;
        ChannelMessage t;
        t <- mod_3151.get(0);
        mod_3150.put(1, t);
    endrule
    rule rule_4074;
        ChannelMessage t;
        t <- mod_3156.get(0);
        mod_3156.put(1, t);
    endrule
    rule rule_4075;
        ChannelMessage t;
        t <- mod_3156.get(1);
        mod_3120.put(1, t);
    endrule
    rule rule_4076;
        ChannelMessage t;
        t <- mod_3127.get(0);
        mod_3128.put(0, t);
    endrule
    rule rule_4077;
        ChannelMessage t;
        t <- mod_3134.get(1);
        mod_3132.put(1, t);
    endrule
    rule rule_4078;
        ChannelMessage t;
        t <- mod_3120.get(1);
        mod_3121.put(0, t);
    endrule
    rule rule_4079;
        ChannelMessage t;
        t <- mod_3135.get(0);
        mod_3135.put(1, t);
    endrule
    rule rule_4080;
        ChannelMessage t;
        t <- mod_3148.get(1);
        mod_3143.put(0, t);
    endrule
    rule rule_4081;
        ChannelMessage t;
        t <- mod_3148.get(0);
        mod_3149.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3117.put(0, t);
        end
        if (i == 1) begin
            mod_3133.put(0, t);
        end
        if (i == 2) begin
            mod_3139.put(0, t);
        end
        if (i == 3) begin
            mod_3147.put(0, t);
        end
        if (i == 4) begin
            mod_3153.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_3121.get(0);
        end
        if (i == 2) begin
            t <- mod_3121.get(1);
        end
        if (i == 0) begin
            t <- mod_3121.get(2);
        end
        if (i == 3) begin
            t <- mod_3133.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6111 (Operation_IFC);
    Operation_IFC mod_3158_inner <- mkReshape(2, 64);
    Operation_IFC mod_3158 <- mkDebugOperation(mod_3158_inner, "mod_3158");
    Operation_IFC mod_3159_inner <- mkFlatten(1);
    Operation_IFC mod_3159 <- mkDebugOperation(mod_3159_inner, "mod_3159");
    Operation_IFC mod_3160_inner <- mkFlatten(2);
    Operation_IFC mod_3160 <- mkDebugOperation(mod_3160_inner, "mod_3160");
    Operation_IFC mod_3161_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3161 <- mkDebugOperation(mod_3161_inner, "mod_3161");
    Broadcast_IFC#(4) mod_3162_inner <- mkBroadcast(4);
    Operation_IFC mod_3162 <- mkDebugOperation(mod_3162_inner.op, "mod_3162");
    PMU_IFC mod_3163_bufferize <- mkPMU(2);
    Operation_IFC mod_3163_inner = mod_3163_bufferize.operation;
    Operation_IFC mod_3163 <- mkDebugOperation(mod_3163_inner, "mod_3163");
    Broadcast_IFC#(2) mod_3164_inner <- mkBroadcast(2);
    Operation_IFC mod_3164 <- mkDebugOperation(mod_3164_inner.op, "mod_3164");
    PMU_IFC mod_3165_bufferize <- mkPMU(1);
    Operation_IFC mod_3165_inner = mod_3165_bufferize.operation;
    Operation_IFC mod_3165 <- mkDebugOperation(mod_3165_inner, "mod_3165");
    Operation_IFC mod_3166_inner <- mkBinaryMap(1079, matmul_t_tile);
    Operation_IFC mod_3166 <- mkDebugOperation(mod_3166_inner, "mod_3166");
    Operation_IFC mod_3167_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3167 <- mkDebugOperation(mod_3167_inner, "mod_3167");
    Operation_IFC mod_3168_inner <- mkBinaryMap(1847, mul_tile);
    Operation_IFC mod_3168 <- mkDebugOperation(mod_3168_inner, "mod_3168");
    PMU_IFC mod_3169_bufferize <- mkPMU(1);
    Operation_IFC mod_3169_inner = mod_3169_bufferize.operation;
    Operation_IFC mod_3169 <- mkDebugOperation(mod_3169_inner, "mod_3169");
    Operation_IFC mod_3170_inner <- mkBinaryMap(2409, matmul_t_tile);
    Operation_IFC mod_3170 <- mkDebugOperation(mod_3170_inner, "mod_3170");
    Operation_IFC mod_3171_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3171 <- mkDebugOperation(mod_3171_inner, "mod_3171");
    Operation_IFC mod_3172_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3172 <- mkDebugOperation(mod_3172_inner, "mod_3172");
    Operation_IFC mod_3173_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3173 <- mkDebugOperation(mod_3173_inner, "mod_3173");
    Operation_IFC mod_3174_inner <- mkBinaryMap(2746, mul_tile);
    Operation_IFC mod_3174 <- mkDebugOperation(mod_3174_inner, "mod_3174");
    PMU_IFC mod_3175_bufferize <- mkPMU(1);
    Operation_IFC mod_3175_inner = mod_3175_bufferize.operation;
    Operation_IFC mod_3175 <- mkDebugOperation(mod_3175_inner, "mod_3175");
    PMU_IFC mod_3176_bufferize <- mkPMU(2);
    Operation_IFC mod_3176_inner = mod_3176_bufferize.operation;
    Operation_IFC mod_3176 <- mkDebugOperation(mod_3176_inner, "mod_3176");
    PMU_IFC mod_3177_bufferize <- mkPMU(2);
    Operation_IFC mod_3177_inner = mod_3177_bufferize.operation;
    Operation_IFC mod_3177 <- mkDebugOperation(mod_3177_inner, "mod_3177");
    Operation_IFC mod_3178_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3178 <- mkDebugOperation(mod_3178_inner, "mod_3178");
    Operation_IFC mod_3179_inner <- mkFlatten(1);
    Operation_IFC mod_3179 <- mkDebugOperation(mod_3179_inner, "mod_3179");
    Operation_IFC mod_3180_inner <- mkFlatten(0);
    Operation_IFC mod_3180 <- mkDebugOperation(mod_3180_inner, "mod_3180");
    Operation_IFC mod_3181_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3181 <- mkDebugOperation(mod_3181_inner, "mod_3181");
    Operation_IFC mod_3182_inner <- mkUnaryMap(1719, silu_tile);
    Operation_IFC mod_3182 <- mkDebugOperation(mod_3182_inner, "mod_3182");
    Operation_IFC mod_3183_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3183 <- mkDebugOperation(mod_3183_inner, "mod_3183");
    Operation_IFC mod_3184_inner <- mkBinaryMap(1591, matmul_t_tile);
    Operation_IFC mod_3184 <- mkDebugOperation(mod_3184_inner, "mod_3184");
    PMU_IFC mod_3185_bufferize <- mkPMU(2);
    Operation_IFC mod_3185_inner = mod_3185_bufferize.operation;
    Operation_IFC mod_3185 <- mkDebugOperation(mod_3185_inner, "mod_3185");
    Operation_IFC mod_3186_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3186 <- mkDebugOperation(mod_3186_inner, "mod_3186");
    Operation_IFC mod_3187_inner <- mkFlatten(1);
    Operation_IFC mod_3187 <- mkDebugOperation(mod_3187_inner, "mod_3187");
    Operation_IFC mod_3188_inner <- mkFlatten(0);
    Operation_IFC mod_3188 <- mkDebugOperation(mod_3188_inner, "mod_3188");
    PMU_IFC mod_3189_bufferize <- mkPMU(1);
    Operation_IFC mod_3189_inner = mod_3189_bufferize.operation;
    Operation_IFC mod_3189 <- mkDebugOperation(mod_3189_inner, "mod_3189");
    Operation_IFC mod_3190_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3190 <- mkDebugOperation(mod_3190_inner, "mod_3190");
    PMU_IFC mod_3191_bufferize <- mkPMU(2);
    Operation_IFC mod_3191_inner = mod_3191_bufferize.operation;
    Operation_IFC mod_3191 <- mkDebugOperation(mod_3191_inner, "mod_3191");
    Operation_IFC mod_3192_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3192 <- mkDebugOperation(mod_3192_inner, "mod_3192");
    Operation_IFC mod_3193_inner <- mkFlatten(1);
    Operation_IFC mod_3193 <- mkDebugOperation(mod_3193_inner, "mod_3193");
    Operation_IFC mod_3194_inner <- mkFlatten(0);
    Operation_IFC mod_3194 <- mkDebugOperation(mod_3194_inner, "mod_3194");
    Operation_IFC mod_3195_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3195 <- mkDebugOperation(mod_3195_inner, "mod_3195");
    Operation_IFC mod_3196_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3196 <- mkDebugOperation(mod_3196_inner, "mod_3196");
    PMU_IFC mod_3197_bufferize <- mkPMU(2);
    Operation_IFC mod_3197_inner = mod_3197_bufferize.operation;
    Operation_IFC mod_3197 <- mkDebugOperation(mod_3197_inner, "mod_3197");
    rule rule_4082;
        ChannelMessage t;
        t <- mod_3175.get(0);
        mod_3175.put(1, t);
    endrule
    rule rule_4083;
        ChannelMessage t;
        t <- mod_3178.get(0);
        mod_3177.put(1, t);
    endrule
    rule rule_4084;
        ChannelMessage t;
        t <- mod_3163.get(0);
        mod_3196.put(0, t);
    endrule
    rule rule_4085;
        ChannelMessage t;
        t <- mod_3165.get(0);
        mod_3195.put(0, t);
    endrule
    rule rule_4086;
        ChannelMessage t;
        t <- mod_3173.get(1);
        mod_3174.put(1, t);
    endrule
    rule rule_4087;
        ChannelMessage t;
        t <- mod_3182.get(0);
        mod_3168.put(1, t);
    endrule
    rule rule_4088;
        ChannelMessage t;
        t <- mod_3165.get(1);
        mod_3166.put(0, t);
    endrule
    rule rule_4089;
        ChannelMessage t;
        t <- mod_3183.get(0);
        mod_3182.put(0, t);
    endrule
    rule rule_4090;
        ChannelMessage t;
        t <- mod_3197.get(0);
        mod_3197.put(1, t);
    endrule
    rule rule_4091;
        ChannelMessage t;
        t <- mod_3177.get(1);
        mod_3170.put(1, t);
    endrule
    rule rule_4092;
        ChannelMessage t;
        t <- mod_3176.get(0);
        mod_3176.put(1, t);
    endrule
    rule rule_4093;
        ChannelMessage t;
        t <- mod_3177.get(0);
        mod_3178.put(0, t);
    endrule
    rule rule_4094;
        ChannelMessage t;
        t <- mod_3186.get(0);
        mod_3185.put(1, t);
    endrule
    rule rule_4095;
        ChannelMessage t;
        t <- mod_3160.get(0);
        mod_3161.put(0, t);
    endrule
    rule rule_4096;
        ChannelMessage t;
        t <- mod_3189.get(0);
        mod_3190.put(0, t);
    endrule
    rule rule_4097;
        ChannelMessage t;
        t <- mod_3190.get(0);
        mod_3189.put(1, t);
    endrule
    rule rule_4098;
        ChannelMessage t;
        t <- mod_3168.get(0);
        mod_3169.put(0, t);
    endrule
    rule rule_4099;
        ChannelMessage t;
        t <- mod_3169.get(1);
        mod_3170.put(0, t);
    endrule
    rule rule_4100;
        ChannelMessage t;
        t <- mod_3159.get(0);
        mod_3160.put(0, t);
    endrule
    rule rule_4101;
        ChannelMessage t;
        t <- mod_3187.get(0);
        mod_3185.put(0, t);
    endrule
    rule rule_4102;
        ChannelMessage t;
        t <- mod_3191.get(0);
        mod_3192.put(0, t);
    endrule
    rule rule_4103;
        ChannelMessage t;
        t <- mod_3185.get(0);
        mod_3186.put(0, t);
    endrule
    rule rule_4104;
        ChannelMessage t;
        t <- mod_3175.get(1);
        mod_3173.put(1, t);
    endrule
    rule rule_4105;
        ChannelMessage t;
        t <- mod_3195.get(0);
        mod_3165.put(1, t);
    endrule
    rule rule_4106;
        ChannelMessage t;
        t <- mod_3188.get(0);
        mod_3187.put(0, t);
    endrule
    rule rule_4107;
        ChannelMessage t;
        t <- mod_3170.get(0);
        mod_3171.put(0, t);
    endrule
    rule rule_4108;
        ChannelMessage t;
        t <- mod_3167.get(0);
        mod_3168.put(0, t);
    endrule
    rule rule_4109;
        ChannelMessage t;
        t <- mod_3180.get(0);
        mod_3179.put(0, t);
    endrule
    rule rule_4110;
        ChannelMessage t;
        t <- mod_3172.get(1);
        mod_3173.put(0, t);
    endrule
    rule rule_4111;
        ChannelMessage t;
        t <- mod_3163.get(1);
        mod_3164.put(0, t);
    endrule
    rule rule_4112;
        ChannelMessage t;
        t <- mod_3181.get(0);
        mod_3169.put(1, t);
    endrule
    rule rule_4113;
        ChannelMessage t;
        t <- mod_3161.get(1);
        mod_3162.put(0, t);
    endrule
    rule rule_4114;
        ChannelMessage t;
        t <- mod_3176.get(1);
        mod_3172.put(1, t);
    endrule
    rule rule_4115;
        ChannelMessage t;
        t <- mod_3197.get(1);
        mod_3161.put(1, t);
    endrule
    rule rule_4116;
        ChannelMessage t;
        t <- mod_3164.get(0);
        mod_3189.put(0, t);
    endrule
    rule rule_4117;
        ChannelMessage t;
        t <- mod_3192.get(0);
        mod_3191.put(1, t);
    endrule
    rule rule_4118;
        ChannelMessage t;
        t <- mod_3179.get(0);
        mod_3177.put(0, t);
    endrule
    rule rule_4119;
        ChannelMessage t;
        t <- mod_3196.get(0);
        mod_3163.put(1, t);
    endrule
    rule rule_4120;
        ChannelMessage t;
        t <- mod_3161.get(0);
        mod_3197.put(0, t);
    endrule
    rule rule_4121;
        ChannelMessage t;
        t <- mod_3171.get(0);
        mod_3172.put(0, t);
    endrule
    rule rule_4122;
        ChannelMessage t;
        t <- mod_3164.get(1);
        mod_3165.put(0, t);
    endrule
    rule rule_4123;
        ChannelMessage t;
        t <- mod_3189.get(1);
        mod_3184.put(0, t);
    endrule
    rule rule_4124;
        ChannelMessage t;
        t <- mod_3162.get(3);
        mod_3163.put(0, t);
    endrule
    rule rule_4125;
        ChannelMessage t;
        t <- mod_3173.get(0);
        mod_3175.put(0, t);
    endrule
    rule rule_4126;
        ChannelMessage t;
        t <- mod_3191.get(1);
        mod_3166.put(1, t);
    endrule
    rule rule_4127;
        ChannelMessage t;
        t <- mod_3158.get(0);
        mod_3159.put(0, t);
    endrule
    rule rule_4128;
        ChannelMessage t;
        t <- mod_3166.get(0);
        mod_3167.put(0, t);
    endrule
    rule rule_4129;
        ChannelMessage t;
        t <- mod_3193.get(0);
        mod_3191.put(0, t);
    endrule
    rule rule_4130;
        ChannelMessage t;
        t <- mod_3169.get(0);
        mod_3181.put(0, t);
    endrule
    rule rule_4131;
        ChannelMessage t;
        t <- mod_3184.get(0);
        mod_3183.put(0, t);
    endrule
    rule rule_4132;
        ChannelMessage t;
        t <- mod_3194.get(0);
        mod_3193.put(0, t);
    endrule
    rule rule_4133;
        ChannelMessage t;
        t <- mod_3185.get(1);
        mod_3184.put(1, t);
    endrule
    rule rule_4134;
        ChannelMessage t;
        t <- mod_3172.get(0);
        mod_3176.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3158.put(0, t);
        end
        if (i == 1) begin
            mod_3174.put(0, t);
        end
        if (i == 2) begin
            mod_3180.put(0, t);
        end
        if (i == 3) begin
            mod_3188.put(0, t);
        end
        if (i == 4) begin
            mod_3194.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_3162.get(0);
        end
        if (i == 1) begin
            t <- mod_3162.get(1);
        end
        if (i == 0) begin
            t <- mod_3162.get(2);
        end
        if (i == 2) begin
            t <- mod_3174.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6112 (Operation_IFC);
    Operation_IFC mod_3199_inner <- mkReshape(2, 64);
    Operation_IFC mod_3199 <- mkDebugOperation(mod_3199_inner, "mod_3199");
    Operation_IFC mod_3200_inner <- mkFlatten(1);
    Operation_IFC mod_3200 <- mkDebugOperation(mod_3200_inner, "mod_3200");
    Operation_IFC mod_3201_inner <- mkFlatten(2);
    Operation_IFC mod_3201 <- mkDebugOperation(mod_3201_inner, "mod_3201");
    Operation_IFC mod_3202_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3202 <- mkDebugOperation(mod_3202_inner, "mod_3202");
    Broadcast_IFC#(4) mod_3203_inner <- mkBroadcast(4);
    Operation_IFC mod_3203 <- mkDebugOperation(mod_3203_inner.op, "mod_3203");
    PMU_IFC mod_3204_bufferize <- mkPMU(2);
    Operation_IFC mod_3204_inner = mod_3204_bufferize.operation;
    Operation_IFC mod_3204 <- mkDebugOperation(mod_3204_inner, "mod_3204");
    Broadcast_IFC#(2) mod_3205_inner <- mkBroadcast(2);
    Operation_IFC mod_3205 <- mkDebugOperation(mod_3205_inner.op, "mod_3205");
    PMU_IFC mod_3206_bufferize <- mkPMU(1);
    Operation_IFC mod_3206_inner = mod_3206_bufferize.operation;
    Operation_IFC mod_3206 <- mkDebugOperation(mod_3206_inner, "mod_3206");
    Operation_IFC mod_3207_inner <- mkBinaryMap(1078, matmul_t_tile);
    Operation_IFC mod_3207 <- mkDebugOperation(mod_3207_inner, "mod_3207");
    Operation_IFC mod_3208_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3208 <- mkDebugOperation(mod_3208_inner, "mod_3208");
    Operation_IFC mod_3209_inner <- mkBinaryMap(1846, mul_tile);
    Operation_IFC mod_3209 <- mkDebugOperation(mod_3209_inner, "mod_3209");
    PMU_IFC mod_3210_bufferize <- mkPMU(1);
    Operation_IFC mod_3210_inner = mod_3210_bufferize.operation;
    Operation_IFC mod_3210 <- mkDebugOperation(mod_3210_inner, "mod_3210");
    Operation_IFC mod_3211_inner <- mkBinaryMap(2407, matmul_t_tile);
    Operation_IFC mod_3211 <- mkDebugOperation(mod_3211_inner, "mod_3211");
    Operation_IFC mod_3212_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3212 <- mkDebugOperation(mod_3212_inner, "mod_3212");
    Operation_IFC mod_3213_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3213 <- mkDebugOperation(mod_3213_inner, "mod_3213");
    Operation_IFC mod_3214_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3214 <- mkDebugOperation(mod_3214_inner, "mod_3214");
    Operation_IFC mod_3215_inner <- mkBinaryMap(2745, mul_tile);
    Operation_IFC mod_3215 <- mkDebugOperation(mod_3215_inner, "mod_3215");
    PMU_IFC mod_3216_bufferize <- mkPMU(1);
    Operation_IFC mod_3216_inner = mod_3216_bufferize.operation;
    Operation_IFC mod_3216 <- mkDebugOperation(mod_3216_inner, "mod_3216");
    PMU_IFC mod_3217_bufferize <- mkPMU(2);
    Operation_IFC mod_3217_inner = mod_3217_bufferize.operation;
    Operation_IFC mod_3217 <- mkDebugOperation(mod_3217_inner, "mod_3217");
    PMU_IFC mod_3218_bufferize <- mkPMU(2);
    Operation_IFC mod_3218_inner = mod_3218_bufferize.operation;
    Operation_IFC mod_3218 <- mkDebugOperation(mod_3218_inner, "mod_3218");
    Operation_IFC mod_3219_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3219 <- mkDebugOperation(mod_3219_inner, "mod_3219");
    Operation_IFC mod_3220_inner <- mkFlatten(1);
    Operation_IFC mod_3220 <- mkDebugOperation(mod_3220_inner, "mod_3220");
    Operation_IFC mod_3221_inner <- mkFlatten(0);
    Operation_IFC mod_3221 <- mkDebugOperation(mod_3221_inner, "mod_3221");
    Operation_IFC mod_3222_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3222 <- mkDebugOperation(mod_3222_inner, "mod_3222");
    Operation_IFC mod_3223_inner <- mkUnaryMap(1718, silu_tile);
    Operation_IFC mod_3223 <- mkDebugOperation(mod_3223_inner, "mod_3223");
    Operation_IFC mod_3224_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3224 <- mkDebugOperation(mod_3224_inner, "mod_3224");
    Operation_IFC mod_3225_inner <- mkBinaryMap(1590, matmul_t_tile);
    Operation_IFC mod_3225 <- mkDebugOperation(mod_3225_inner, "mod_3225");
    PMU_IFC mod_3226_bufferize <- mkPMU(2);
    Operation_IFC mod_3226_inner = mod_3226_bufferize.operation;
    Operation_IFC mod_3226 <- mkDebugOperation(mod_3226_inner, "mod_3226");
    Operation_IFC mod_3227_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3227 <- mkDebugOperation(mod_3227_inner, "mod_3227");
    Operation_IFC mod_3228_inner <- mkFlatten(1);
    Operation_IFC mod_3228 <- mkDebugOperation(mod_3228_inner, "mod_3228");
    Operation_IFC mod_3229_inner <- mkFlatten(0);
    Operation_IFC mod_3229 <- mkDebugOperation(mod_3229_inner, "mod_3229");
    PMU_IFC mod_3230_bufferize <- mkPMU(1);
    Operation_IFC mod_3230_inner = mod_3230_bufferize.operation;
    Operation_IFC mod_3230 <- mkDebugOperation(mod_3230_inner, "mod_3230");
    Operation_IFC mod_3231_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3231 <- mkDebugOperation(mod_3231_inner, "mod_3231");
    PMU_IFC mod_3232_bufferize <- mkPMU(2);
    Operation_IFC mod_3232_inner = mod_3232_bufferize.operation;
    Operation_IFC mod_3232 <- mkDebugOperation(mod_3232_inner, "mod_3232");
    Operation_IFC mod_3233_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3233 <- mkDebugOperation(mod_3233_inner, "mod_3233");
    Operation_IFC mod_3234_inner <- mkFlatten(1);
    Operation_IFC mod_3234 <- mkDebugOperation(mod_3234_inner, "mod_3234");
    Operation_IFC mod_3235_inner <- mkFlatten(0);
    Operation_IFC mod_3235 <- mkDebugOperation(mod_3235_inner, "mod_3235");
    Operation_IFC mod_3236_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3236 <- mkDebugOperation(mod_3236_inner, "mod_3236");
    Operation_IFC mod_3237_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3237 <- mkDebugOperation(mod_3237_inner, "mod_3237");
    PMU_IFC mod_3238_bufferize <- mkPMU(2);
    Operation_IFC mod_3238_inner = mod_3238_bufferize.operation;
    Operation_IFC mod_3238 <- mkDebugOperation(mod_3238_inner, "mod_3238");
    rule rule_4135;
        ChannelMessage t;
        t <- mod_3205.get(1);
        mod_3206.put(0, t);
    endrule
    rule rule_4136;
        ChannelMessage t;
        t <- mod_3217.get(1);
        mod_3213.put(1, t);
    endrule
    rule rule_4137;
        ChannelMessage t;
        t <- mod_3211.get(0);
        mod_3212.put(0, t);
    endrule
    rule rule_4138;
        ChannelMessage t;
        t <- mod_3218.get(0);
        mod_3219.put(0, t);
    endrule
    rule rule_4139;
        ChannelMessage t;
        t <- mod_3226.get(1);
        mod_3225.put(1, t);
    endrule
    rule rule_4140;
        ChannelMessage t;
        t <- mod_3214.get(0);
        mod_3216.put(0, t);
    endrule
    rule rule_4141;
        ChannelMessage t;
        t <- mod_3206.get(0);
        mod_3236.put(0, t);
    endrule
    rule rule_4142;
        ChannelMessage t;
        t <- mod_3204.get(0);
        mod_3237.put(0, t);
    endrule
    rule rule_4143;
        ChannelMessage t;
        t <- mod_3216.get(1);
        mod_3214.put(1, t);
    endrule
    rule rule_4144;
        ChannelMessage t;
        t <- mod_3231.get(0);
        mod_3230.put(1, t);
    endrule
    rule rule_4145;
        ChannelMessage t;
        t <- mod_3204.get(1);
        mod_3205.put(0, t);
    endrule
    rule rule_4146;
        ChannelMessage t;
        t <- mod_3212.get(0);
        mod_3213.put(0, t);
    endrule
    rule rule_4147;
        ChannelMessage t;
        t <- mod_3222.get(0);
        mod_3210.put(1, t);
    endrule
    rule rule_4148;
        ChannelMessage t;
        t <- mod_3232.get(1);
        mod_3207.put(1, t);
    endrule
    rule rule_4149;
        ChannelMessage t;
        t <- mod_3202.get(1);
        mod_3203.put(0, t);
    endrule
    rule rule_4150;
        ChannelMessage t;
        t <- mod_3221.get(0);
        mod_3220.put(0, t);
    endrule
    rule rule_4151;
        ChannelMessage t;
        t <- mod_3205.get(0);
        mod_3230.put(0, t);
    endrule
    rule rule_4152;
        ChannelMessage t;
        t <- mod_3214.get(1);
        mod_3215.put(1, t);
    endrule
    rule rule_4153;
        ChannelMessage t;
        t <- mod_3225.get(0);
        mod_3224.put(0, t);
    endrule
    rule rule_4154;
        ChannelMessage t;
        t <- mod_3208.get(0);
        mod_3209.put(0, t);
    endrule
    rule rule_4155;
        ChannelMessage t;
        t <- mod_3210.get(0);
        mod_3222.put(0, t);
    endrule
    rule rule_4156;
        ChannelMessage t;
        t <- mod_3213.get(0);
        mod_3217.put(0, t);
    endrule
    rule rule_4157;
        ChannelMessage t;
        t <- mod_3200.get(0);
        mod_3201.put(0, t);
    endrule
    rule rule_4158;
        ChannelMessage t;
        t <- mod_3228.get(0);
        mod_3226.put(0, t);
    endrule
    rule rule_4159;
        ChannelMessage t;
        t <- mod_3233.get(0);
        mod_3232.put(1, t);
    endrule
    rule rule_4160;
        ChannelMessage t;
        t <- mod_3219.get(0);
        mod_3218.put(1, t);
    endrule
    rule rule_4161;
        ChannelMessage t;
        t <- mod_3224.get(0);
        mod_3223.put(0, t);
    endrule
    rule rule_4162;
        ChannelMessage t;
        t <- mod_3227.get(0);
        mod_3226.put(1, t);
    endrule
    rule rule_4163;
        ChannelMessage t;
        t <- mod_3217.get(0);
        mod_3217.put(1, t);
    endrule
    rule rule_4164;
        ChannelMessage t;
        t <- mod_3220.get(0);
        mod_3218.put(0, t);
    endrule
    rule rule_4165;
        ChannelMessage t;
        t <- mod_3238.get(0);
        mod_3238.put(1, t);
    endrule
    rule rule_4166;
        ChannelMessage t;
        t <- mod_3199.get(0);
        mod_3200.put(0, t);
    endrule
    rule rule_4167;
        ChannelMessage t;
        t <- mod_3229.get(0);
        mod_3228.put(0, t);
    endrule
    rule rule_4168;
        ChannelMessage t;
        t <- mod_3206.get(1);
        mod_3207.put(0, t);
    endrule
    rule rule_4169;
        ChannelMessage t;
        t <- mod_3216.get(0);
        mod_3216.put(1, t);
    endrule
    rule rule_4170;
        ChannelMessage t;
        t <- mod_3237.get(0);
        mod_3204.put(1, t);
    endrule
    rule rule_4171;
        ChannelMessage t;
        t <- mod_3234.get(0);
        mod_3232.put(0, t);
    endrule
    rule rule_4172;
        ChannelMessage t;
        t <- mod_3202.get(0);
        mod_3238.put(0, t);
    endrule
    rule rule_4173;
        ChannelMessage t;
        t <- mod_3213.get(1);
        mod_3214.put(0, t);
    endrule
    rule rule_4174;
        ChannelMessage t;
        t <- mod_3235.get(0);
        mod_3234.put(0, t);
    endrule
    rule rule_4175;
        ChannelMessage t;
        t <- mod_3210.get(1);
        mod_3211.put(0, t);
    endrule
    rule rule_4176;
        ChannelMessage t;
        t <- mod_3201.get(0);
        mod_3202.put(0, t);
    endrule
    rule rule_4177;
        ChannelMessage t;
        t <- mod_3223.get(0);
        mod_3209.put(1, t);
    endrule
    rule rule_4178;
        ChannelMessage t;
        t <- mod_3207.get(0);
        mod_3208.put(0, t);
    endrule
    rule rule_4179;
        ChannelMessage t;
        t <- mod_3226.get(0);
        mod_3227.put(0, t);
    endrule
    rule rule_4180;
        ChannelMessage t;
        t <- mod_3232.get(0);
        mod_3233.put(0, t);
    endrule
    rule rule_4181;
        ChannelMessage t;
        t <- mod_3230.get(0);
        mod_3231.put(0, t);
    endrule
    rule rule_4182;
        ChannelMessage t;
        t <- mod_3236.get(0);
        mod_3206.put(1, t);
    endrule
    rule rule_4183;
        ChannelMessage t;
        t <- mod_3209.get(0);
        mod_3210.put(0, t);
    endrule
    rule rule_4184;
        ChannelMessage t;
        t <- mod_3203.get(3);
        mod_3204.put(0, t);
    endrule
    rule rule_4185;
        ChannelMessage t;
        t <- mod_3238.get(1);
        mod_3202.put(1, t);
    endrule
    rule rule_4186;
        ChannelMessage t;
        t <- mod_3230.get(1);
        mod_3225.put(0, t);
    endrule
    rule rule_4187;
        ChannelMessage t;
        t <- mod_3218.get(1);
        mod_3211.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3199.put(0, t);
        end
        if (i == 1) begin
            mod_3215.put(0, t);
        end
        if (i == 2) begin
            mod_3221.put(0, t);
        end
        if (i == 3) begin
            mod_3229.put(0, t);
        end
        if (i == 4) begin
            mod_3235.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_3203.get(0);
        end
        if (i == 0) begin
            t <- mod_3203.get(1);
        end
        if (i == 3) begin
            t <- mod_3203.get(2);
        end
        if (i == 2) begin
            t <- mod_3215.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6113 (Operation_IFC);
    Operation_IFC mod_3240_inner <- mkReshape(2, 64);
    Operation_IFC mod_3240 <- mkDebugOperation(mod_3240_inner, "mod_3240");
    Operation_IFC mod_3241_inner <- mkFlatten(1);
    Operation_IFC mod_3241 <- mkDebugOperation(mod_3241_inner, "mod_3241");
    Operation_IFC mod_3242_inner <- mkFlatten(2);
    Operation_IFC mod_3242 <- mkDebugOperation(mod_3242_inner, "mod_3242");
    Operation_IFC mod_3243_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3243 <- mkDebugOperation(mod_3243_inner, "mod_3243");
    Broadcast_IFC#(4) mod_3244_inner <- mkBroadcast(4);
    Operation_IFC mod_3244 <- mkDebugOperation(mod_3244_inner.op, "mod_3244");
    PMU_IFC mod_3245_bufferize <- mkPMU(2);
    Operation_IFC mod_3245_inner = mod_3245_bufferize.operation;
    Operation_IFC mod_3245 <- mkDebugOperation(mod_3245_inner, "mod_3245");
    Broadcast_IFC#(2) mod_3246_inner <- mkBroadcast(2);
    Operation_IFC mod_3246 <- mkDebugOperation(mod_3246_inner.op, "mod_3246");
    PMU_IFC mod_3247_bufferize <- mkPMU(1);
    Operation_IFC mod_3247_inner = mod_3247_bufferize.operation;
    Operation_IFC mod_3247 <- mkDebugOperation(mod_3247_inner, "mod_3247");
    Operation_IFC mod_3248_inner <- mkBinaryMap(1077, matmul_t_tile);
    Operation_IFC mod_3248 <- mkDebugOperation(mod_3248_inner, "mod_3248");
    Operation_IFC mod_3249_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3249 <- mkDebugOperation(mod_3249_inner, "mod_3249");
    Operation_IFC mod_3250_inner <- mkBinaryMap(1845, mul_tile);
    Operation_IFC mod_3250 <- mkDebugOperation(mod_3250_inner, "mod_3250");
    PMU_IFC mod_3251_bufferize <- mkPMU(1);
    Operation_IFC mod_3251_inner = mod_3251_bufferize.operation;
    Operation_IFC mod_3251 <- mkDebugOperation(mod_3251_inner, "mod_3251");
    Operation_IFC mod_3252_inner <- mkBinaryMap(2405, matmul_t_tile);
    Operation_IFC mod_3252 <- mkDebugOperation(mod_3252_inner, "mod_3252");
    Operation_IFC mod_3253_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3253 <- mkDebugOperation(mod_3253_inner, "mod_3253");
    Operation_IFC mod_3254_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3254 <- mkDebugOperation(mod_3254_inner, "mod_3254");
    Operation_IFC mod_3255_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3255 <- mkDebugOperation(mod_3255_inner, "mod_3255");
    Operation_IFC mod_3256_inner <- mkBinaryMap(2744, mul_tile);
    Operation_IFC mod_3256 <- mkDebugOperation(mod_3256_inner, "mod_3256");
    PMU_IFC mod_3257_bufferize <- mkPMU(1);
    Operation_IFC mod_3257_inner = mod_3257_bufferize.operation;
    Operation_IFC mod_3257 <- mkDebugOperation(mod_3257_inner, "mod_3257");
    PMU_IFC mod_3258_bufferize <- mkPMU(2);
    Operation_IFC mod_3258_inner = mod_3258_bufferize.operation;
    Operation_IFC mod_3258 <- mkDebugOperation(mod_3258_inner, "mod_3258");
    PMU_IFC mod_3259_bufferize <- mkPMU(2);
    Operation_IFC mod_3259_inner = mod_3259_bufferize.operation;
    Operation_IFC mod_3259 <- mkDebugOperation(mod_3259_inner, "mod_3259");
    Operation_IFC mod_3260_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3260 <- mkDebugOperation(mod_3260_inner, "mod_3260");
    Operation_IFC mod_3261_inner <- mkFlatten(1);
    Operation_IFC mod_3261 <- mkDebugOperation(mod_3261_inner, "mod_3261");
    Operation_IFC mod_3262_inner <- mkFlatten(0);
    Operation_IFC mod_3262 <- mkDebugOperation(mod_3262_inner, "mod_3262");
    Operation_IFC mod_3263_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3263 <- mkDebugOperation(mod_3263_inner, "mod_3263");
    Operation_IFC mod_3264_inner <- mkUnaryMap(1717, silu_tile);
    Operation_IFC mod_3264 <- mkDebugOperation(mod_3264_inner, "mod_3264");
    Operation_IFC mod_3265_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3265 <- mkDebugOperation(mod_3265_inner, "mod_3265");
    Operation_IFC mod_3266_inner <- mkBinaryMap(1589, matmul_t_tile);
    Operation_IFC mod_3266 <- mkDebugOperation(mod_3266_inner, "mod_3266");
    PMU_IFC mod_3267_bufferize <- mkPMU(2);
    Operation_IFC mod_3267_inner = mod_3267_bufferize.operation;
    Operation_IFC mod_3267 <- mkDebugOperation(mod_3267_inner, "mod_3267");
    Operation_IFC mod_3268_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3268 <- mkDebugOperation(mod_3268_inner, "mod_3268");
    Operation_IFC mod_3269_inner <- mkFlatten(1);
    Operation_IFC mod_3269 <- mkDebugOperation(mod_3269_inner, "mod_3269");
    Operation_IFC mod_3270_inner <- mkFlatten(0);
    Operation_IFC mod_3270 <- mkDebugOperation(mod_3270_inner, "mod_3270");
    PMU_IFC mod_3271_bufferize <- mkPMU(1);
    Operation_IFC mod_3271_inner = mod_3271_bufferize.operation;
    Operation_IFC mod_3271 <- mkDebugOperation(mod_3271_inner, "mod_3271");
    Operation_IFC mod_3272_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3272 <- mkDebugOperation(mod_3272_inner, "mod_3272");
    PMU_IFC mod_3273_bufferize <- mkPMU(2);
    Operation_IFC mod_3273_inner = mod_3273_bufferize.operation;
    Operation_IFC mod_3273 <- mkDebugOperation(mod_3273_inner, "mod_3273");
    Operation_IFC mod_3274_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3274 <- mkDebugOperation(mod_3274_inner, "mod_3274");
    Operation_IFC mod_3275_inner <- mkFlatten(1);
    Operation_IFC mod_3275 <- mkDebugOperation(mod_3275_inner, "mod_3275");
    Operation_IFC mod_3276_inner <- mkFlatten(0);
    Operation_IFC mod_3276 <- mkDebugOperation(mod_3276_inner, "mod_3276");
    Operation_IFC mod_3277_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3277 <- mkDebugOperation(mod_3277_inner, "mod_3277");
    Operation_IFC mod_3278_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3278 <- mkDebugOperation(mod_3278_inner, "mod_3278");
    PMU_IFC mod_3279_bufferize <- mkPMU(2);
    Operation_IFC mod_3279_inner = mod_3279_bufferize.operation;
    Operation_IFC mod_3279 <- mkDebugOperation(mod_3279_inner, "mod_3279");
    rule rule_4188;
        ChannelMessage t;
        t <- mod_3240.get(0);
        mod_3241.put(0, t);
    endrule
    rule rule_4189;
        ChannelMessage t;
        t <- mod_3279.get(1);
        mod_3243.put(1, t);
    endrule
    rule rule_4190;
        ChannelMessage t;
        t <- mod_3252.get(0);
        mod_3253.put(0, t);
    endrule
    rule rule_4191;
        ChannelMessage t;
        t <- mod_3265.get(0);
        mod_3264.put(0, t);
    endrule
    rule rule_4192;
        ChannelMessage t;
        t <- mod_3251.get(0);
        mod_3263.put(0, t);
    endrule
    rule rule_4193;
        ChannelMessage t;
        t <- mod_3250.get(0);
        mod_3251.put(0, t);
    endrule
    rule rule_4194;
        ChannelMessage t;
        t <- mod_3251.get(1);
        mod_3252.put(0, t);
    endrule
    rule rule_4195;
        ChannelMessage t;
        t <- mod_3255.get(1);
        mod_3256.put(1, t);
    endrule
    rule rule_4196;
        ChannelMessage t;
        t <- mod_3267.get(1);
        mod_3266.put(1, t);
    endrule
    rule rule_4197;
        ChannelMessage t;
        t <- mod_3254.get(0);
        mod_3258.put(0, t);
    endrule
    rule rule_4198;
        ChannelMessage t;
        t <- mod_3245.get(0);
        mod_3278.put(0, t);
    endrule
    rule rule_4199;
        ChannelMessage t;
        t <- mod_3259.get(1);
        mod_3252.put(1, t);
    endrule
    rule rule_4200;
        ChannelMessage t;
        t <- mod_3248.get(0);
        mod_3249.put(0, t);
    endrule
    rule rule_4201;
        ChannelMessage t;
        t <- mod_3255.get(0);
        mod_3257.put(0, t);
    endrule
    rule rule_4202;
        ChannelMessage t;
        t <- mod_3243.get(0);
        mod_3279.put(0, t);
    endrule
    rule rule_4203;
        ChannelMessage t;
        t <- mod_3241.get(0);
        mod_3242.put(0, t);
    endrule
    rule rule_4204;
        ChannelMessage t;
        t <- mod_3247.get(1);
        mod_3248.put(0, t);
    endrule
    rule rule_4205;
        ChannelMessage t;
        t <- mod_3266.get(0);
        mod_3265.put(0, t);
    endrule
    rule rule_4206;
        ChannelMessage t;
        t <- mod_3277.get(0);
        mod_3247.put(1, t);
    endrule
    rule rule_4207;
        ChannelMessage t;
        t <- mod_3270.get(0);
        mod_3269.put(0, t);
    endrule
    rule rule_4208;
        ChannelMessage t;
        t <- mod_3279.get(0);
        mod_3279.put(1, t);
    endrule
    rule rule_4209;
        ChannelMessage t;
        t <- mod_3242.get(0);
        mod_3243.put(0, t);
    endrule
    rule rule_4210;
        ChannelMessage t;
        t <- mod_3267.get(0);
        mod_3268.put(0, t);
    endrule
    rule rule_4211;
        ChannelMessage t;
        t <- mod_3276.get(0);
        mod_3275.put(0, t);
    endrule
    rule rule_4212;
        ChannelMessage t;
        t <- mod_3247.get(0);
        mod_3277.put(0, t);
    endrule
    rule rule_4213;
        ChannelMessage t;
        t <- mod_3245.get(1);
        mod_3246.put(0, t);
    endrule
    rule rule_4214;
        ChannelMessage t;
        t <- mod_3275.get(0);
        mod_3273.put(0, t);
    endrule
    rule rule_4215;
        ChannelMessage t;
        t <- mod_3246.get(1);
        mod_3247.put(0, t);
    endrule
    rule rule_4216;
        ChannelMessage t;
        t <- mod_3254.get(1);
        mod_3255.put(0, t);
    endrule
    rule rule_4217;
        ChannelMessage t;
        t <- mod_3258.get(0);
        mod_3258.put(1, t);
    endrule
    rule rule_4218;
        ChannelMessage t;
        t <- mod_3274.get(0);
        mod_3273.put(1, t);
    endrule
    rule rule_4219;
        ChannelMessage t;
        t <- mod_3246.get(0);
        mod_3271.put(0, t);
    endrule
    rule rule_4220;
        ChannelMessage t;
        t <- mod_3258.get(1);
        mod_3254.put(1, t);
    endrule
    rule rule_4221;
        ChannelMessage t;
        t <- mod_3278.get(0);
        mod_3245.put(1, t);
    endrule
    rule rule_4222;
        ChannelMessage t;
        t <- mod_3263.get(0);
        mod_3251.put(1, t);
    endrule
    rule rule_4223;
        ChannelMessage t;
        t <- mod_3244.get(3);
        mod_3245.put(0, t);
    endrule
    rule rule_4224;
        ChannelMessage t;
        t <- mod_3249.get(0);
        mod_3250.put(0, t);
    endrule
    rule rule_4225;
        ChannelMessage t;
        t <- mod_3264.get(0);
        mod_3250.put(1, t);
    endrule
    rule rule_4226;
        ChannelMessage t;
        t <- mod_3271.get(1);
        mod_3266.put(0, t);
    endrule
    rule rule_4227;
        ChannelMessage t;
        t <- mod_3272.get(0);
        mod_3271.put(1, t);
    endrule
    rule rule_4228;
        ChannelMessage t;
        t <- mod_3243.get(1);
        mod_3244.put(0, t);
    endrule
    rule rule_4229;
        ChannelMessage t;
        t <- mod_3257.get(0);
        mod_3257.put(1, t);
    endrule
    rule rule_4230;
        ChannelMessage t;
        t <- mod_3253.get(0);
        mod_3254.put(0, t);
    endrule
    rule rule_4231;
        ChannelMessage t;
        t <- mod_3261.get(0);
        mod_3259.put(0, t);
    endrule
    rule rule_4232;
        ChannelMessage t;
        t <- mod_3273.get(0);
        mod_3274.put(0, t);
    endrule
    rule rule_4233;
        ChannelMessage t;
        t <- mod_3257.get(1);
        mod_3255.put(1, t);
    endrule
    rule rule_4234;
        ChannelMessage t;
        t <- mod_3260.get(0);
        mod_3259.put(1, t);
    endrule
    rule rule_4235;
        ChannelMessage t;
        t <- mod_3269.get(0);
        mod_3267.put(0, t);
    endrule
    rule rule_4236;
        ChannelMessage t;
        t <- mod_3271.get(0);
        mod_3272.put(0, t);
    endrule
    rule rule_4237;
        ChannelMessage t;
        t <- mod_3262.get(0);
        mod_3261.put(0, t);
    endrule
    rule rule_4238;
        ChannelMessage t;
        t <- mod_3259.get(0);
        mod_3260.put(0, t);
    endrule
    rule rule_4239;
        ChannelMessage t;
        t <- mod_3268.get(0);
        mod_3267.put(1, t);
    endrule
    rule rule_4240;
        ChannelMessage t;
        t <- mod_3273.get(1);
        mod_3248.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3240.put(0, t);
        end
        if (i == 1) begin
            mod_3256.put(0, t);
        end
        if (i == 2) begin
            mod_3262.put(0, t);
        end
        if (i == 3) begin
            mod_3270.put(0, t);
        end
        if (i == 4) begin
            mod_3276.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_3244.get(0);
        end
        if (i == 0) begin
            t <- mod_3244.get(1);
        end
        if (i == 1) begin
            t <- mod_3244.get(2);
        end
        if (i == 2) begin
            t <- mod_3256.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6114 (Operation_IFC);
    Operation_IFC mod_3281_inner <- mkReshape(2, 64);
    Operation_IFC mod_3281 <- mkDebugOperation(mod_3281_inner, "mod_3281");
    Operation_IFC mod_3282_inner <- mkFlatten(1);
    Operation_IFC mod_3282 <- mkDebugOperation(mod_3282_inner, "mod_3282");
    Operation_IFC mod_3283_inner <- mkFlatten(2);
    Operation_IFC mod_3283 <- mkDebugOperation(mod_3283_inner, "mod_3283");
    Operation_IFC mod_3284_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3284 <- mkDebugOperation(mod_3284_inner, "mod_3284");
    Broadcast_IFC#(4) mod_3285_inner <- mkBroadcast(4);
    Operation_IFC mod_3285 <- mkDebugOperation(mod_3285_inner.op, "mod_3285");
    PMU_IFC mod_3286_bufferize <- mkPMU(2);
    Operation_IFC mod_3286_inner = mod_3286_bufferize.operation;
    Operation_IFC mod_3286 <- mkDebugOperation(mod_3286_inner, "mod_3286");
    Broadcast_IFC#(2) mod_3287_inner <- mkBroadcast(2);
    Operation_IFC mod_3287 <- mkDebugOperation(mod_3287_inner.op, "mod_3287");
    PMU_IFC mod_3288_bufferize <- mkPMU(1);
    Operation_IFC mod_3288_inner = mod_3288_bufferize.operation;
    Operation_IFC mod_3288 <- mkDebugOperation(mod_3288_inner, "mod_3288");
    Operation_IFC mod_3289_inner <- mkBinaryMap(1076, matmul_t_tile);
    Operation_IFC mod_3289 <- mkDebugOperation(mod_3289_inner, "mod_3289");
    Operation_IFC mod_3290_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3290 <- mkDebugOperation(mod_3290_inner, "mod_3290");
    Operation_IFC mod_3291_inner <- mkBinaryMap(1844, mul_tile);
    Operation_IFC mod_3291 <- mkDebugOperation(mod_3291_inner, "mod_3291");
    PMU_IFC mod_3292_bufferize <- mkPMU(1);
    Operation_IFC mod_3292_inner = mod_3292_bufferize.operation;
    Operation_IFC mod_3292 <- mkDebugOperation(mod_3292_inner, "mod_3292");
    Operation_IFC mod_3293_inner <- mkBinaryMap(2403, matmul_t_tile);
    Operation_IFC mod_3293 <- mkDebugOperation(mod_3293_inner, "mod_3293");
    Operation_IFC mod_3294_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3294 <- mkDebugOperation(mod_3294_inner, "mod_3294");
    Operation_IFC mod_3295_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3295 <- mkDebugOperation(mod_3295_inner, "mod_3295");
    Operation_IFC mod_3296_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3296 <- mkDebugOperation(mod_3296_inner, "mod_3296");
    Operation_IFC mod_3297_inner <- mkBinaryMap(2743, mul_tile);
    Operation_IFC mod_3297 <- mkDebugOperation(mod_3297_inner, "mod_3297");
    PMU_IFC mod_3298_bufferize <- mkPMU(1);
    Operation_IFC mod_3298_inner = mod_3298_bufferize.operation;
    Operation_IFC mod_3298 <- mkDebugOperation(mod_3298_inner, "mod_3298");
    PMU_IFC mod_3299_bufferize <- mkPMU(2);
    Operation_IFC mod_3299_inner = mod_3299_bufferize.operation;
    Operation_IFC mod_3299 <- mkDebugOperation(mod_3299_inner, "mod_3299");
    PMU_IFC mod_3300_bufferize <- mkPMU(2);
    Operation_IFC mod_3300_inner = mod_3300_bufferize.operation;
    Operation_IFC mod_3300 <- mkDebugOperation(mod_3300_inner, "mod_3300");
    Operation_IFC mod_3301_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3301 <- mkDebugOperation(mod_3301_inner, "mod_3301");
    Operation_IFC mod_3302_inner <- mkFlatten(1);
    Operation_IFC mod_3302 <- mkDebugOperation(mod_3302_inner, "mod_3302");
    Operation_IFC mod_3303_inner <- mkFlatten(0);
    Operation_IFC mod_3303 <- mkDebugOperation(mod_3303_inner, "mod_3303");
    Operation_IFC mod_3304_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3304 <- mkDebugOperation(mod_3304_inner, "mod_3304");
    Operation_IFC mod_3305_inner <- mkUnaryMap(1716, silu_tile);
    Operation_IFC mod_3305 <- mkDebugOperation(mod_3305_inner, "mod_3305");
    Operation_IFC mod_3306_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3306 <- mkDebugOperation(mod_3306_inner, "mod_3306");
    Operation_IFC mod_3307_inner <- mkBinaryMap(1588, matmul_t_tile);
    Operation_IFC mod_3307 <- mkDebugOperation(mod_3307_inner, "mod_3307");
    PMU_IFC mod_3308_bufferize <- mkPMU(2);
    Operation_IFC mod_3308_inner = mod_3308_bufferize.operation;
    Operation_IFC mod_3308 <- mkDebugOperation(mod_3308_inner, "mod_3308");
    Operation_IFC mod_3309_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3309 <- mkDebugOperation(mod_3309_inner, "mod_3309");
    Operation_IFC mod_3310_inner <- mkFlatten(1);
    Operation_IFC mod_3310 <- mkDebugOperation(mod_3310_inner, "mod_3310");
    Operation_IFC mod_3311_inner <- mkFlatten(0);
    Operation_IFC mod_3311 <- mkDebugOperation(mod_3311_inner, "mod_3311");
    PMU_IFC mod_3312_bufferize <- mkPMU(1);
    Operation_IFC mod_3312_inner = mod_3312_bufferize.operation;
    Operation_IFC mod_3312 <- mkDebugOperation(mod_3312_inner, "mod_3312");
    Operation_IFC mod_3313_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3313 <- mkDebugOperation(mod_3313_inner, "mod_3313");
    PMU_IFC mod_3314_bufferize <- mkPMU(2);
    Operation_IFC mod_3314_inner = mod_3314_bufferize.operation;
    Operation_IFC mod_3314 <- mkDebugOperation(mod_3314_inner, "mod_3314");
    Operation_IFC mod_3315_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3315 <- mkDebugOperation(mod_3315_inner, "mod_3315");
    Operation_IFC mod_3316_inner <- mkFlatten(1);
    Operation_IFC mod_3316 <- mkDebugOperation(mod_3316_inner, "mod_3316");
    Operation_IFC mod_3317_inner <- mkFlatten(0);
    Operation_IFC mod_3317 <- mkDebugOperation(mod_3317_inner, "mod_3317");
    Operation_IFC mod_3318_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3318 <- mkDebugOperation(mod_3318_inner, "mod_3318");
    Operation_IFC mod_3319_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3319 <- mkDebugOperation(mod_3319_inner, "mod_3319");
    PMU_IFC mod_3320_bufferize <- mkPMU(2);
    Operation_IFC mod_3320_inner = mod_3320_bufferize.operation;
    Operation_IFC mod_3320 <- mkDebugOperation(mod_3320_inner, "mod_3320");
    rule rule_4241;
        ChannelMessage t;
        t <- mod_3288.get(0);
        mod_3318.put(0, t);
    endrule
    rule rule_4242;
        ChannelMessage t;
        t <- mod_3300.get(0);
        mod_3301.put(0, t);
    endrule
    rule rule_4243;
        ChannelMessage t;
        t <- mod_3291.get(0);
        mod_3292.put(0, t);
    endrule
    rule rule_4244;
        ChannelMessage t;
        t <- mod_3284.get(0);
        mod_3320.put(0, t);
    endrule
    rule rule_4245;
        ChannelMessage t;
        t <- mod_3296.get(0);
        mod_3298.put(0, t);
    endrule
    rule rule_4246;
        ChannelMessage t;
        t <- mod_3312.get(0);
        mod_3313.put(0, t);
    endrule
    rule rule_4247;
        ChannelMessage t;
        t <- mod_3282.get(0);
        mod_3283.put(0, t);
    endrule
    rule rule_4248;
        ChannelMessage t;
        t <- mod_3289.get(0);
        mod_3290.put(0, t);
    endrule
    rule rule_4249;
        ChannelMessage t;
        t <- mod_3300.get(1);
        mod_3293.put(1, t);
    endrule
    rule rule_4250;
        ChannelMessage t;
        t <- mod_3302.get(0);
        mod_3300.put(0, t);
    endrule
    rule rule_4251;
        ChannelMessage t;
        t <- mod_3308.get(0);
        mod_3309.put(0, t);
    endrule
    rule rule_4252;
        ChannelMessage t;
        t <- mod_3311.get(0);
        mod_3310.put(0, t);
    endrule
    rule rule_4253;
        ChannelMessage t;
        t <- mod_3318.get(0);
        mod_3288.put(1, t);
    endrule
    rule rule_4254;
        ChannelMessage t;
        t <- mod_3319.get(0);
        mod_3286.put(1, t);
    endrule
    rule rule_4255;
        ChannelMessage t;
        t <- mod_3283.get(0);
        mod_3284.put(0, t);
    endrule
    rule rule_4256;
        ChannelMessage t;
        t <- mod_3309.get(0);
        mod_3308.put(1, t);
    endrule
    rule rule_4257;
        ChannelMessage t;
        t <- mod_3295.get(0);
        mod_3299.put(0, t);
    endrule
    rule rule_4258;
        ChannelMessage t;
        t <- mod_3298.get(1);
        mod_3296.put(1, t);
    endrule
    rule rule_4259;
        ChannelMessage t;
        t <- mod_3288.get(1);
        mod_3289.put(0, t);
    endrule
    rule rule_4260;
        ChannelMessage t;
        t <- mod_3296.get(1);
        mod_3297.put(1, t);
    endrule
    rule rule_4261;
        ChannelMessage t;
        t <- mod_3287.get(0);
        mod_3312.put(0, t);
    endrule
    rule rule_4262;
        ChannelMessage t;
        t <- mod_3313.get(0);
        mod_3312.put(1, t);
    endrule
    rule rule_4263;
        ChannelMessage t;
        t <- mod_3286.get(1);
        mod_3287.put(0, t);
    endrule
    rule rule_4264;
        ChannelMessage t;
        t <- mod_3299.get(0);
        mod_3299.put(1, t);
    endrule
    rule rule_4265;
        ChannelMessage t;
        t <- mod_3299.get(1);
        mod_3295.put(1, t);
    endrule
    rule rule_4266;
        ChannelMessage t;
        t <- mod_3314.get(0);
        mod_3315.put(0, t);
    endrule
    rule rule_4267;
        ChannelMessage t;
        t <- mod_3294.get(0);
        mod_3295.put(0, t);
    endrule
    rule rule_4268;
        ChannelMessage t;
        t <- mod_3320.get(1);
        mod_3284.put(1, t);
    endrule
    rule rule_4269;
        ChannelMessage t;
        t <- mod_3301.get(0);
        mod_3300.put(1, t);
    endrule
    rule rule_4270;
        ChannelMessage t;
        t <- mod_3293.get(0);
        mod_3294.put(0, t);
    endrule
    rule rule_4271;
        ChannelMessage t;
        t <- mod_3316.get(0);
        mod_3314.put(0, t);
    endrule
    rule rule_4272;
        ChannelMessage t;
        t <- mod_3304.get(0);
        mod_3292.put(1, t);
    endrule
    rule rule_4273;
        ChannelMessage t;
        t <- mod_3310.get(0);
        mod_3308.put(0, t);
    endrule
    rule rule_4274;
        ChannelMessage t;
        t <- mod_3298.get(0);
        mod_3298.put(1, t);
    endrule
    rule rule_4275;
        ChannelMessage t;
        t <- mod_3286.get(0);
        mod_3319.put(0, t);
    endrule
    rule rule_4276;
        ChannelMessage t;
        t <- mod_3290.get(0);
        mod_3291.put(0, t);
    endrule
    rule rule_4277;
        ChannelMessage t;
        t <- mod_3285.get(3);
        mod_3286.put(0, t);
    endrule
    rule rule_4278;
        ChannelMessage t;
        t <- mod_3292.get(0);
        mod_3304.put(0, t);
    endrule
    rule rule_4279;
        ChannelMessage t;
        t <- mod_3314.get(1);
        mod_3289.put(1, t);
    endrule
    rule rule_4280;
        ChannelMessage t;
        t <- mod_3317.get(0);
        mod_3316.put(0, t);
    endrule
    rule rule_4281;
        ChannelMessage t;
        t <- mod_3284.get(1);
        mod_3285.put(0, t);
    endrule
    rule rule_4282;
        ChannelMessage t;
        t <- mod_3281.get(0);
        mod_3282.put(0, t);
    endrule
    rule rule_4283;
        ChannelMessage t;
        t <- mod_3307.get(0);
        mod_3306.put(0, t);
    endrule
    rule rule_4284;
        ChannelMessage t;
        t <- mod_3305.get(0);
        mod_3291.put(1, t);
    endrule
    rule rule_4285;
        ChannelMessage t;
        t <- mod_3312.get(1);
        mod_3307.put(0, t);
    endrule
    rule rule_4286;
        ChannelMessage t;
        t <- mod_3315.get(0);
        mod_3314.put(1, t);
    endrule
    rule rule_4287;
        ChannelMessage t;
        t <- mod_3303.get(0);
        mod_3302.put(0, t);
    endrule
    rule rule_4288;
        ChannelMessage t;
        t <- mod_3292.get(1);
        mod_3293.put(0, t);
    endrule
    rule rule_4289;
        ChannelMessage t;
        t <- mod_3287.get(1);
        mod_3288.put(0, t);
    endrule
    rule rule_4290;
        ChannelMessage t;
        t <- mod_3295.get(1);
        mod_3296.put(0, t);
    endrule
    rule rule_4291;
        ChannelMessage t;
        t <- mod_3308.get(1);
        mod_3307.put(1, t);
    endrule
    rule rule_4292;
        ChannelMessage t;
        t <- mod_3320.get(0);
        mod_3320.put(1, t);
    endrule
    rule rule_4293;
        ChannelMessage t;
        t <- mod_3306.get(0);
        mod_3305.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3281.put(0, t);
        end
        if (i == 1) begin
            mod_3297.put(0, t);
        end
        if (i == 2) begin
            mod_3303.put(0, t);
        end
        if (i == 3) begin
            mod_3311.put(0, t);
        end
        if (i == 4) begin
            mod_3317.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_3285.get(0);
        end
        if (i == 2) begin
            t <- mod_3285.get(1);
        end
        if (i == 0) begin
            t <- mod_3285.get(2);
        end
        if (i == 3) begin
            t <- mod_3297.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6115 (Operation_IFC);
    Operation_IFC mod_3322_inner <- mkReshape(2, 64);
    Operation_IFC mod_3322 <- mkDebugOperation(mod_3322_inner, "mod_3322");
    Operation_IFC mod_3323_inner <- mkFlatten(1);
    Operation_IFC mod_3323 <- mkDebugOperation(mod_3323_inner, "mod_3323");
    Operation_IFC mod_3324_inner <- mkFlatten(2);
    Operation_IFC mod_3324 <- mkDebugOperation(mod_3324_inner, "mod_3324");
    Operation_IFC mod_3325_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3325 <- mkDebugOperation(mod_3325_inner, "mod_3325");
    Broadcast_IFC#(4) mod_3326_inner <- mkBroadcast(4);
    Operation_IFC mod_3326 <- mkDebugOperation(mod_3326_inner.op, "mod_3326");
    PMU_IFC mod_3327_bufferize <- mkPMU(2);
    Operation_IFC mod_3327_inner = mod_3327_bufferize.operation;
    Operation_IFC mod_3327 <- mkDebugOperation(mod_3327_inner, "mod_3327");
    Broadcast_IFC#(2) mod_3328_inner <- mkBroadcast(2);
    Operation_IFC mod_3328 <- mkDebugOperation(mod_3328_inner.op, "mod_3328");
    PMU_IFC mod_3329_bufferize <- mkPMU(1);
    Operation_IFC mod_3329_inner = mod_3329_bufferize.operation;
    Operation_IFC mod_3329 <- mkDebugOperation(mod_3329_inner, "mod_3329");
    Operation_IFC mod_3330_inner <- mkBinaryMap(1075, matmul_t_tile);
    Operation_IFC mod_3330 <- mkDebugOperation(mod_3330_inner, "mod_3330");
    Operation_IFC mod_3331_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3331 <- mkDebugOperation(mod_3331_inner, "mod_3331");
    Operation_IFC mod_3332_inner <- mkBinaryMap(1843, mul_tile);
    Operation_IFC mod_3332 <- mkDebugOperation(mod_3332_inner, "mod_3332");
    PMU_IFC mod_3333_bufferize <- mkPMU(1);
    Operation_IFC mod_3333_inner = mod_3333_bufferize.operation;
    Operation_IFC mod_3333 <- mkDebugOperation(mod_3333_inner, "mod_3333");
    Operation_IFC mod_3334_inner <- mkBinaryMap(2401, matmul_t_tile);
    Operation_IFC mod_3334 <- mkDebugOperation(mod_3334_inner, "mod_3334");
    Operation_IFC mod_3335_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3335 <- mkDebugOperation(mod_3335_inner, "mod_3335");
    Operation_IFC mod_3336_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3336 <- mkDebugOperation(mod_3336_inner, "mod_3336");
    Operation_IFC mod_3337_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3337 <- mkDebugOperation(mod_3337_inner, "mod_3337");
    Operation_IFC mod_3338_inner <- mkBinaryMap(2742, mul_tile);
    Operation_IFC mod_3338 <- mkDebugOperation(mod_3338_inner, "mod_3338");
    PMU_IFC mod_3339_bufferize <- mkPMU(1);
    Operation_IFC mod_3339_inner = mod_3339_bufferize.operation;
    Operation_IFC mod_3339 <- mkDebugOperation(mod_3339_inner, "mod_3339");
    PMU_IFC mod_3340_bufferize <- mkPMU(2);
    Operation_IFC mod_3340_inner = mod_3340_bufferize.operation;
    Operation_IFC mod_3340 <- mkDebugOperation(mod_3340_inner, "mod_3340");
    PMU_IFC mod_3341_bufferize <- mkPMU(2);
    Operation_IFC mod_3341_inner = mod_3341_bufferize.operation;
    Operation_IFC mod_3341 <- mkDebugOperation(mod_3341_inner, "mod_3341");
    Operation_IFC mod_3342_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3342 <- mkDebugOperation(mod_3342_inner, "mod_3342");
    Operation_IFC mod_3343_inner <- mkFlatten(1);
    Operation_IFC mod_3343 <- mkDebugOperation(mod_3343_inner, "mod_3343");
    Operation_IFC mod_3344_inner <- mkFlatten(0);
    Operation_IFC mod_3344 <- mkDebugOperation(mod_3344_inner, "mod_3344");
    Operation_IFC mod_3345_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3345 <- mkDebugOperation(mod_3345_inner, "mod_3345");
    Operation_IFC mod_3346_inner <- mkUnaryMap(1715, silu_tile);
    Operation_IFC mod_3346 <- mkDebugOperation(mod_3346_inner, "mod_3346");
    Operation_IFC mod_3347_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3347 <- mkDebugOperation(mod_3347_inner, "mod_3347");
    Operation_IFC mod_3348_inner <- mkBinaryMap(1587, matmul_t_tile);
    Operation_IFC mod_3348 <- mkDebugOperation(mod_3348_inner, "mod_3348");
    PMU_IFC mod_3349_bufferize <- mkPMU(2);
    Operation_IFC mod_3349_inner = mod_3349_bufferize.operation;
    Operation_IFC mod_3349 <- mkDebugOperation(mod_3349_inner, "mod_3349");
    Operation_IFC mod_3350_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3350 <- mkDebugOperation(mod_3350_inner, "mod_3350");
    Operation_IFC mod_3351_inner <- mkFlatten(1);
    Operation_IFC mod_3351 <- mkDebugOperation(mod_3351_inner, "mod_3351");
    Operation_IFC mod_3352_inner <- mkFlatten(0);
    Operation_IFC mod_3352 <- mkDebugOperation(mod_3352_inner, "mod_3352");
    PMU_IFC mod_3353_bufferize <- mkPMU(1);
    Operation_IFC mod_3353_inner = mod_3353_bufferize.operation;
    Operation_IFC mod_3353 <- mkDebugOperation(mod_3353_inner, "mod_3353");
    Operation_IFC mod_3354_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3354 <- mkDebugOperation(mod_3354_inner, "mod_3354");
    PMU_IFC mod_3355_bufferize <- mkPMU(2);
    Operation_IFC mod_3355_inner = mod_3355_bufferize.operation;
    Operation_IFC mod_3355 <- mkDebugOperation(mod_3355_inner, "mod_3355");
    Operation_IFC mod_3356_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3356 <- mkDebugOperation(mod_3356_inner, "mod_3356");
    Operation_IFC mod_3357_inner <- mkFlatten(1);
    Operation_IFC mod_3357 <- mkDebugOperation(mod_3357_inner, "mod_3357");
    Operation_IFC mod_3358_inner <- mkFlatten(0);
    Operation_IFC mod_3358 <- mkDebugOperation(mod_3358_inner, "mod_3358");
    Operation_IFC mod_3359_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3359 <- mkDebugOperation(mod_3359_inner, "mod_3359");
    Operation_IFC mod_3360_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3360 <- mkDebugOperation(mod_3360_inner, "mod_3360");
    PMU_IFC mod_3361_bufferize <- mkPMU(2);
    Operation_IFC mod_3361_inner = mod_3361_bufferize.operation;
    Operation_IFC mod_3361 <- mkDebugOperation(mod_3361_inner, "mod_3361");
    rule rule_4294;
        ChannelMessage t;
        t <- mod_3331.get(0);
        mod_3332.put(0, t);
    endrule
    rule rule_4295;
        ChannelMessage t;
        t <- mod_3323.get(0);
        mod_3324.put(0, t);
    endrule
    rule rule_4296;
        ChannelMessage t;
        t <- mod_3361.get(0);
        mod_3361.put(1, t);
    endrule
    rule rule_4297;
        ChannelMessage t;
        t <- mod_3346.get(0);
        mod_3332.put(1, t);
    endrule
    rule rule_4298;
        ChannelMessage t;
        t <- mod_3328.get(1);
        mod_3329.put(0, t);
    endrule
    rule rule_4299;
        ChannelMessage t;
        t <- mod_3349.get(1);
        mod_3348.put(1, t);
    endrule
    rule rule_4300;
        ChannelMessage t;
        t <- mod_3333.get(0);
        mod_3345.put(0, t);
    endrule
    rule rule_4301;
        ChannelMessage t;
        t <- mod_3356.get(0);
        mod_3355.put(1, t);
    endrule
    rule rule_4302;
        ChannelMessage t;
        t <- mod_3352.get(0);
        mod_3351.put(0, t);
    endrule
    rule rule_4303;
        ChannelMessage t;
        t <- mod_3361.get(1);
        mod_3325.put(1, t);
    endrule
    rule rule_4304;
        ChannelMessage t;
        t <- mod_3333.get(1);
        mod_3334.put(0, t);
    endrule
    rule rule_4305;
        ChannelMessage t;
        t <- mod_3355.get(0);
        mod_3356.put(0, t);
    endrule
    rule rule_4306;
        ChannelMessage t;
        t <- mod_3330.get(0);
        mod_3331.put(0, t);
    endrule
    rule rule_4307;
        ChannelMessage t;
        t <- mod_3350.get(0);
        mod_3349.put(1, t);
    endrule
    rule rule_4308;
        ChannelMessage t;
        t <- mod_3340.get(1);
        mod_3336.put(1, t);
    endrule
    rule rule_4309;
        ChannelMessage t;
        t <- mod_3327.get(1);
        mod_3328.put(0, t);
    endrule
    rule rule_4310;
        ChannelMessage t;
        t <- mod_3339.get(1);
        mod_3337.put(1, t);
    endrule
    rule rule_4311;
        ChannelMessage t;
        t <- mod_3325.get(0);
        mod_3361.put(0, t);
    endrule
    rule rule_4312;
        ChannelMessage t;
        t <- mod_3345.get(0);
        mod_3333.put(1, t);
    endrule
    rule rule_4313;
        ChannelMessage t;
        t <- mod_3347.get(0);
        mod_3346.put(0, t);
    endrule
    rule rule_4314;
        ChannelMessage t;
        t <- mod_3357.get(0);
        mod_3355.put(0, t);
    endrule
    rule rule_4315;
        ChannelMessage t;
        t <- mod_3325.get(1);
        mod_3326.put(0, t);
    endrule
    rule rule_4316;
        ChannelMessage t;
        t <- mod_3344.get(0);
        mod_3343.put(0, t);
    endrule
    rule rule_4317;
        ChannelMessage t;
        t <- mod_3359.get(0);
        mod_3329.put(1, t);
    endrule
    rule rule_4318;
        ChannelMessage t;
        t <- mod_3342.get(0);
        mod_3341.put(1, t);
    endrule
    rule rule_4319;
        ChannelMessage t;
        t <- mod_3336.get(0);
        mod_3340.put(0, t);
    endrule
    rule rule_4320;
        ChannelMessage t;
        t <- mod_3336.get(1);
        mod_3337.put(0, t);
    endrule
    rule rule_4321;
        ChannelMessage t;
        t <- mod_3341.get(0);
        mod_3342.put(0, t);
    endrule
    rule rule_4322;
        ChannelMessage t;
        t <- mod_3353.get(1);
        mod_3348.put(0, t);
    endrule
    rule rule_4323;
        ChannelMessage t;
        t <- mod_3360.get(0);
        mod_3327.put(1, t);
    endrule
    rule rule_4324;
        ChannelMessage t;
        t <- mod_3348.get(0);
        mod_3347.put(0, t);
    endrule
    rule rule_4325;
        ChannelMessage t;
        t <- mod_3349.get(0);
        mod_3350.put(0, t);
    endrule
    rule rule_4326;
        ChannelMessage t;
        t <- mod_3355.get(1);
        mod_3330.put(1, t);
    endrule
    rule rule_4327;
        ChannelMessage t;
        t <- mod_3335.get(0);
        mod_3336.put(0, t);
    endrule
    rule rule_4328;
        ChannelMessage t;
        t <- mod_3327.get(0);
        mod_3360.put(0, t);
    endrule
    rule rule_4329;
        ChannelMessage t;
        t <- mod_3324.get(0);
        mod_3325.put(0, t);
    endrule
    rule rule_4330;
        ChannelMessage t;
        t <- mod_3339.get(0);
        mod_3339.put(1, t);
    endrule
    rule rule_4331;
        ChannelMessage t;
        t <- mod_3332.get(0);
        mod_3333.put(0, t);
    endrule
    rule rule_4332;
        ChannelMessage t;
        t <- mod_3337.get(0);
        mod_3339.put(0, t);
    endrule
    rule rule_4333;
        ChannelMessage t;
        t <- mod_3341.get(1);
        mod_3334.put(1, t);
    endrule
    rule rule_4334;
        ChannelMessage t;
        t <- mod_3353.get(0);
        mod_3354.put(0, t);
    endrule
    rule rule_4335;
        ChannelMessage t;
        t <- mod_3329.get(0);
        mod_3359.put(0, t);
    endrule
    rule rule_4336;
        ChannelMessage t;
        t <- mod_3322.get(0);
        mod_3323.put(0, t);
    endrule
    rule rule_4337;
        ChannelMessage t;
        t <- mod_3358.get(0);
        mod_3357.put(0, t);
    endrule
    rule rule_4338;
        ChannelMessage t;
        t <- mod_3340.get(0);
        mod_3340.put(1, t);
    endrule
    rule rule_4339;
        ChannelMessage t;
        t <- mod_3337.get(1);
        mod_3338.put(1, t);
    endrule
    rule rule_4340;
        ChannelMessage t;
        t <- mod_3328.get(0);
        mod_3353.put(0, t);
    endrule
    rule rule_4341;
        ChannelMessage t;
        t <- mod_3334.get(0);
        mod_3335.put(0, t);
    endrule
    rule rule_4342;
        ChannelMessage t;
        t <- mod_3326.get(3);
        mod_3327.put(0, t);
    endrule
    rule rule_4343;
        ChannelMessage t;
        t <- mod_3343.get(0);
        mod_3341.put(0, t);
    endrule
    rule rule_4344;
        ChannelMessage t;
        t <- mod_3354.get(0);
        mod_3353.put(1, t);
    endrule
    rule rule_4345;
        ChannelMessage t;
        t <- mod_3329.get(1);
        mod_3330.put(0, t);
    endrule
    rule rule_4346;
        ChannelMessage t;
        t <- mod_3351.get(0);
        mod_3349.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3322.put(0, t);
        end
        if (i == 1) begin
            mod_3338.put(0, t);
        end
        if (i == 2) begin
            mod_3344.put(0, t);
        end
        if (i == 3) begin
            mod_3352.put(0, t);
        end
        if (i == 4) begin
            mod_3358.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_3326.get(0);
        end
        if (i == 2) begin
            t <- mod_3326.get(1);
        end
        if (i == 0) begin
            t <- mod_3326.get(2);
        end
        if (i == 3) begin
            t <- mod_3338.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6116 (Operation_IFC);
    Operation_IFC mod_3363_inner <- mkReshape(2, 64);
    Operation_IFC mod_3363 <- mkDebugOperation(mod_3363_inner, "mod_3363");
    Operation_IFC mod_3364_inner <- mkFlatten(1);
    Operation_IFC mod_3364 <- mkDebugOperation(mod_3364_inner, "mod_3364");
    Operation_IFC mod_3365_inner <- mkFlatten(2);
    Operation_IFC mod_3365 <- mkDebugOperation(mod_3365_inner, "mod_3365");
    Operation_IFC mod_3366_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3366 <- mkDebugOperation(mod_3366_inner, "mod_3366");
    Broadcast_IFC#(4) mod_3367_inner <- mkBroadcast(4);
    Operation_IFC mod_3367 <- mkDebugOperation(mod_3367_inner.op, "mod_3367");
    PMU_IFC mod_3368_bufferize <- mkPMU(2);
    Operation_IFC mod_3368_inner = mod_3368_bufferize.operation;
    Operation_IFC mod_3368 <- mkDebugOperation(mod_3368_inner, "mod_3368");
    Broadcast_IFC#(2) mod_3369_inner <- mkBroadcast(2);
    Operation_IFC mod_3369 <- mkDebugOperation(mod_3369_inner.op, "mod_3369");
    PMU_IFC mod_3370_bufferize <- mkPMU(1);
    Operation_IFC mod_3370_inner = mod_3370_bufferize.operation;
    Operation_IFC mod_3370 <- mkDebugOperation(mod_3370_inner, "mod_3370");
    Operation_IFC mod_3371_inner <- mkBinaryMap(1074, matmul_t_tile);
    Operation_IFC mod_3371 <- mkDebugOperation(mod_3371_inner, "mod_3371");
    Operation_IFC mod_3372_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3372 <- mkDebugOperation(mod_3372_inner, "mod_3372");
    Operation_IFC mod_3373_inner <- mkBinaryMap(1842, mul_tile);
    Operation_IFC mod_3373 <- mkDebugOperation(mod_3373_inner, "mod_3373");
    PMU_IFC mod_3374_bufferize <- mkPMU(1);
    Operation_IFC mod_3374_inner = mod_3374_bufferize.operation;
    Operation_IFC mod_3374 <- mkDebugOperation(mod_3374_inner, "mod_3374");
    Operation_IFC mod_3375_inner <- mkBinaryMap(2399, matmul_t_tile);
    Operation_IFC mod_3375 <- mkDebugOperation(mod_3375_inner, "mod_3375");
    Operation_IFC mod_3376_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3376 <- mkDebugOperation(mod_3376_inner, "mod_3376");
    Operation_IFC mod_3377_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3377 <- mkDebugOperation(mod_3377_inner, "mod_3377");
    Operation_IFC mod_3378_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3378 <- mkDebugOperation(mod_3378_inner, "mod_3378");
    Operation_IFC mod_3379_inner <- mkBinaryMap(2741, mul_tile);
    Operation_IFC mod_3379 <- mkDebugOperation(mod_3379_inner, "mod_3379");
    PMU_IFC mod_3380_bufferize <- mkPMU(1);
    Operation_IFC mod_3380_inner = mod_3380_bufferize.operation;
    Operation_IFC mod_3380 <- mkDebugOperation(mod_3380_inner, "mod_3380");
    PMU_IFC mod_3381_bufferize <- mkPMU(2);
    Operation_IFC mod_3381_inner = mod_3381_bufferize.operation;
    Operation_IFC mod_3381 <- mkDebugOperation(mod_3381_inner, "mod_3381");
    PMU_IFC mod_3382_bufferize <- mkPMU(2);
    Operation_IFC mod_3382_inner = mod_3382_bufferize.operation;
    Operation_IFC mod_3382 <- mkDebugOperation(mod_3382_inner, "mod_3382");
    Operation_IFC mod_3383_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3383 <- mkDebugOperation(mod_3383_inner, "mod_3383");
    Operation_IFC mod_3384_inner <- mkFlatten(1);
    Operation_IFC mod_3384 <- mkDebugOperation(mod_3384_inner, "mod_3384");
    Operation_IFC mod_3385_inner <- mkFlatten(0);
    Operation_IFC mod_3385 <- mkDebugOperation(mod_3385_inner, "mod_3385");
    Operation_IFC mod_3386_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3386 <- mkDebugOperation(mod_3386_inner, "mod_3386");
    Operation_IFC mod_3387_inner <- mkUnaryMap(1714, silu_tile);
    Operation_IFC mod_3387 <- mkDebugOperation(mod_3387_inner, "mod_3387");
    Operation_IFC mod_3388_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3388 <- mkDebugOperation(mod_3388_inner, "mod_3388");
    Operation_IFC mod_3389_inner <- mkBinaryMap(1586, matmul_t_tile);
    Operation_IFC mod_3389 <- mkDebugOperation(mod_3389_inner, "mod_3389");
    PMU_IFC mod_3390_bufferize <- mkPMU(2);
    Operation_IFC mod_3390_inner = mod_3390_bufferize.operation;
    Operation_IFC mod_3390 <- mkDebugOperation(mod_3390_inner, "mod_3390");
    Operation_IFC mod_3391_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3391 <- mkDebugOperation(mod_3391_inner, "mod_3391");
    Operation_IFC mod_3392_inner <- mkFlatten(1);
    Operation_IFC mod_3392 <- mkDebugOperation(mod_3392_inner, "mod_3392");
    Operation_IFC mod_3393_inner <- mkFlatten(0);
    Operation_IFC mod_3393 <- mkDebugOperation(mod_3393_inner, "mod_3393");
    PMU_IFC mod_3394_bufferize <- mkPMU(1);
    Operation_IFC mod_3394_inner = mod_3394_bufferize.operation;
    Operation_IFC mod_3394 <- mkDebugOperation(mod_3394_inner, "mod_3394");
    Operation_IFC mod_3395_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3395 <- mkDebugOperation(mod_3395_inner, "mod_3395");
    PMU_IFC mod_3396_bufferize <- mkPMU(2);
    Operation_IFC mod_3396_inner = mod_3396_bufferize.operation;
    Operation_IFC mod_3396 <- mkDebugOperation(mod_3396_inner, "mod_3396");
    Operation_IFC mod_3397_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3397 <- mkDebugOperation(mod_3397_inner, "mod_3397");
    Operation_IFC mod_3398_inner <- mkFlatten(1);
    Operation_IFC mod_3398 <- mkDebugOperation(mod_3398_inner, "mod_3398");
    Operation_IFC mod_3399_inner <- mkFlatten(0);
    Operation_IFC mod_3399 <- mkDebugOperation(mod_3399_inner, "mod_3399");
    Operation_IFC mod_3400_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3400 <- mkDebugOperation(mod_3400_inner, "mod_3400");
    Operation_IFC mod_3401_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3401 <- mkDebugOperation(mod_3401_inner, "mod_3401");
    PMU_IFC mod_3402_bufferize <- mkPMU(2);
    Operation_IFC mod_3402_inner = mod_3402_bufferize.operation;
    Operation_IFC mod_3402 <- mkDebugOperation(mod_3402_inner, "mod_3402");
    rule rule_4347;
        ChannelMessage t;
        t <- mod_3370.get(1);
        mod_3371.put(0, t);
    endrule
    rule rule_4348;
        ChannelMessage t;
        t <- mod_3390.get(1);
        mod_3389.put(1, t);
    endrule
    rule rule_4349;
        ChannelMessage t;
        t <- mod_3380.get(1);
        mod_3378.put(1, t);
    endrule
    rule rule_4350;
        ChannelMessage t;
        t <- mod_3380.get(0);
        mod_3380.put(1, t);
    endrule
    rule rule_4351;
        ChannelMessage t;
        t <- mod_3367.get(3);
        mod_3368.put(0, t);
    endrule
    rule rule_4352;
        ChannelMessage t;
        t <- mod_3394.get(0);
        mod_3395.put(0, t);
    endrule
    rule rule_4353;
        ChannelMessage t;
        t <- mod_3369.get(0);
        mod_3394.put(0, t);
    endrule
    rule rule_4354;
        ChannelMessage t;
        t <- mod_3386.get(0);
        mod_3374.put(1, t);
    endrule
    rule rule_4355;
        ChannelMessage t;
        t <- mod_3400.get(0);
        mod_3370.put(1, t);
    endrule
    rule rule_4356;
        ChannelMessage t;
        t <- mod_3376.get(0);
        mod_3377.put(0, t);
    endrule
    rule rule_4357;
        ChannelMessage t;
        t <- mod_3382.get(1);
        mod_3375.put(1, t);
    endrule
    rule rule_4358;
        ChannelMessage t;
        t <- mod_3395.get(0);
        mod_3394.put(1, t);
    endrule
    rule rule_4359;
        ChannelMessage t;
        t <- mod_3372.get(0);
        mod_3373.put(0, t);
    endrule
    rule rule_4360;
        ChannelMessage t;
        t <- mod_3363.get(0);
        mod_3364.put(0, t);
    endrule
    rule rule_4361;
        ChannelMessage t;
        t <- mod_3396.get(1);
        mod_3371.put(1, t);
    endrule
    rule rule_4362;
        ChannelMessage t;
        t <- mod_3396.get(0);
        mod_3397.put(0, t);
    endrule
    rule rule_4363;
        ChannelMessage t;
        t <- mod_3381.get(0);
        mod_3381.put(1, t);
    endrule
    rule rule_4364;
        ChannelMessage t;
        t <- mod_3374.get(0);
        mod_3386.put(0, t);
    endrule
    rule rule_4365;
        ChannelMessage t;
        t <- mod_3383.get(0);
        mod_3382.put(1, t);
    endrule
    rule rule_4366;
        ChannelMessage t;
        t <- mod_3402.get(1);
        mod_3366.put(1, t);
    endrule
    rule rule_4367;
        ChannelMessage t;
        t <- mod_3394.get(1);
        mod_3389.put(0, t);
    endrule
    rule rule_4368;
        ChannelMessage t;
        t <- mod_3399.get(0);
        mod_3398.put(0, t);
    endrule
    rule rule_4369;
        ChannelMessage t;
        t <- mod_3370.get(0);
        mod_3400.put(0, t);
    endrule
    rule rule_4370;
        ChannelMessage t;
        t <- mod_3402.get(0);
        mod_3402.put(1, t);
    endrule
    rule rule_4371;
        ChannelMessage t;
        t <- mod_3371.get(0);
        mod_3372.put(0, t);
    endrule
    rule rule_4372;
        ChannelMessage t;
        t <- mod_3377.get(0);
        mod_3381.put(0, t);
    endrule
    rule rule_4373;
        ChannelMessage t;
        t <- mod_3381.get(1);
        mod_3377.put(1, t);
    endrule
    rule rule_4374;
        ChannelMessage t;
        t <- mod_3369.get(1);
        mod_3370.put(0, t);
    endrule
    rule rule_4375;
        ChannelMessage t;
        t <- mod_3382.get(0);
        mod_3383.put(0, t);
    endrule
    rule rule_4376;
        ChannelMessage t;
        t <- mod_3389.get(0);
        mod_3388.put(0, t);
    endrule
    rule rule_4377;
        ChannelMessage t;
        t <- mod_3390.get(0);
        mod_3391.put(0, t);
    endrule
    rule rule_4378;
        ChannelMessage t;
        t <- mod_3392.get(0);
        mod_3390.put(0, t);
    endrule
    rule rule_4379;
        ChannelMessage t;
        t <- mod_3387.get(0);
        mod_3373.put(1, t);
    endrule
    rule rule_4380;
        ChannelMessage t;
        t <- mod_3374.get(1);
        mod_3375.put(0, t);
    endrule
    rule rule_4381;
        ChannelMessage t;
        t <- mod_3385.get(0);
        mod_3384.put(0, t);
    endrule
    rule rule_4382;
        ChannelMessage t;
        t <- mod_3388.get(0);
        mod_3387.put(0, t);
    endrule
    rule rule_4383;
        ChannelMessage t;
        t <- mod_3398.get(0);
        mod_3396.put(0, t);
    endrule
    rule rule_4384;
        ChannelMessage t;
        t <- mod_3378.get(1);
        mod_3379.put(1, t);
    endrule
    rule rule_4385;
        ChannelMessage t;
        t <- mod_3368.get(1);
        mod_3369.put(0, t);
    endrule
    rule rule_4386;
        ChannelMessage t;
        t <- mod_3366.get(0);
        mod_3402.put(0, t);
    endrule
    rule rule_4387;
        ChannelMessage t;
        t <- mod_3375.get(0);
        mod_3376.put(0, t);
    endrule
    rule rule_4388;
        ChannelMessage t;
        t <- mod_3365.get(0);
        mod_3366.put(0, t);
    endrule
    rule rule_4389;
        ChannelMessage t;
        t <- mod_3378.get(0);
        mod_3380.put(0, t);
    endrule
    rule rule_4390;
        ChannelMessage t;
        t <- mod_3393.get(0);
        mod_3392.put(0, t);
    endrule
    rule rule_4391;
        ChannelMessage t;
        t <- mod_3384.get(0);
        mod_3382.put(0, t);
    endrule
    rule rule_4392;
        ChannelMessage t;
        t <- mod_3364.get(0);
        mod_3365.put(0, t);
    endrule
    rule rule_4393;
        ChannelMessage t;
        t <- mod_3366.get(1);
        mod_3367.put(0, t);
    endrule
    rule rule_4394;
        ChannelMessage t;
        t <- mod_3401.get(0);
        mod_3368.put(1, t);
    endrule
    rule rule_4395;
        ChannelMessage t;
        t <- mod_3377.get(1);
        mod_3378.put(0, t);
    endrule
    rule rule_4396;
        ChannelMessage t;
        t <- mod_3391.get(0);
        mod_3390.put(1, t);
    endrule
    rule rule_4397;
        ChannelMessage t;
        t <- mod_3397.get(0);
        mod_3396.put(1, t);
    endrule
    rule rule_4398;
        ChannelMessage t;
        t <- mod_3373.get(0);
        mod_3374.put(0, t);
    endrule
    rule rule_4399;
        ChannelMessage t;
        t <- mod_3368.get(0);
        mod_3401.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3363.put(0, t);
        end
        if (i == 1) begin
            mod_3379.put(0, t);
        end
        if (i == 2) begin
            mod_3385.put(0, t);
        end
        if (i == 3) begin
            mod_3393.put(0, t);
        end
        if (i == 4) begin
            mod_3399.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_3367.get(0);
        end
        if (i == 2) begin
            t <- mod_3367.get(1);
        end
        if (i == 1) begin
            t <- mod_3367.get(2);
        end
        if (i == 0) begin
            t <- mod_3379.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6117 (Operation_IFC);
    Operation_IFC mod_3404_inner <- mkReshape(2, 64);
    Operation_IFC mod_3404 <- mkDebugOperation(mod_3404_inner, "mod_3404");
    Operation_IFC mod_3405_inner <- mkFlatten(1);
    Operation_IFC mod_3405 <- mkDebugOperation(mod_3405_inner, "mod_3405");
    Operation_IFC mod_3406_inner <- mkFlatten(2);
    Operation_IFC mod_3406 <- mkDebugOperation(mod_3406_inner, "mod_3406");
    Operation_IFC mod_3407_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3407 <- mkDebugOperation(mod_3407_inner, "mod_3407");
    Broadcast_IFC#(4) mod_3408_inner <- mkBroadcast(4);
    Operation_IFC mod_3408 <- mkDebugOperation(mod_3408_inner.op, "mod_3408");
    PMU_IFC mod_3409_bufferize <- mkPMU(2);
    Operation_IFC mod_3409_inner = mod_3409_bufferize.operation;
    Operation_IFC mod_3409 <- mkDebugOperation(mod_3409_inner, "mod_3409");
    Broadcast_IFC#(2) mod_3410_inner <- mkBroadcast(2);
    Operation_IFC mod_3410 <- mkDebugOperation(mod_3410_inner.op, "mod_3410");
    PMU_IFC mod_3411_bufferize <- mkPMU(1);
    Operation_IFC mod_3411_inner = mod_3411_bufferize.operation;
    Operation_IFC mod_3411 <- mkDebugOperation(mod_3411_inner, "mod_3411");
    Operation_IFC mod_3412_inner <- mkBinaryMap(1073, matmul_t_tile);
    Operation_IFC mod_3412 <- mkDebugOperation(mod_3412_inner, "mod_3412");
    Operation_IFC mod_3413_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3413 <- mkDebugOperation(mod_3413_inner, "mod_3413");
    Operation_IFC mod_3414_inner <- mkBinaryMap(1841, mul_tile);
    Operation_IFC mod_3414 <- mkDebugOperation(mod_3414_inner, "mod_3414");
    PMU_IFC mod_3415_bufferize <- mkPMU(1);
    Operation_IFC mod_3415_inner = mod_3415_bufferize.operation;
    Operation_IFC mod_3415 <- mkDebugOperation(mod_3415_inner, "mod_3415");
    Operation_IFC mod_3416_inner <- mkBinaryMap(2397, matmul_t_tile);
    Operation_IFC mod_3416 <- mkDebugOperation(mod_3416_inner, "mod_3416");
    Operation_IFC mod_3417_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3417 <- mkDebugOperation(mod_3417_inner, "mod_3417");
    Operation_IFC mod_3418_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3418 <- mkDebugOperation(mod_3418_inner, "mod_3418");
    Operation_IFC mod_3419_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3419 <- mkDebugOperation(mod_3419_inner, "mod_3419");
    Operation_IFC mod_3420_inner <- mkBinaryMap(2740, mul_tile);
    Operation_IFC mod_3420 <- mkDebugOperation(mod_3420_inner, "mod_3420");
    PMU_IFC mod_3421_bufferize <- mkPMU(1);
    Operation_IFC mod_3421_inner = mod_3421_bufferize.operation;
    Operation_IFC mod_3421 <- mkDebugOperation(mod_3421_inner, "mod_3421");
    PMU_IFC mod_3422_bufferize <- mkPMU(2);
    Operation_IFC mod_3422_inner = mod_3422_bufferize.operation;
    Operation_IFC mod_3422 <- mkDebugOperation(mod_3422_inner, "mod_3422");
    PMU_IFC mod_3423_bufferize <- mkPMU(2);
    Operation_IFC mod_3423_inner = mod_3423_bufferize.operation;
    Operation_IFC mod_3423 <- mkDebugOperation(mod_3423_inner, "mod_3423");
    Operation_IFC mod_3424_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3424 <- mkDebugOperation(mod_3424_inner, "mod_3424");
    Operation_IFC mod_3425_inner <- mkFlatten(1);
    Operation_IFC mod_3425 <- mkDebugOperation(mod_3425_inner, "mod_3425");
    Operation_IFC mod_3426_inner <- mkFlatten(0);
    Operation_IFC mod_3426 <- mkDebugOperation(mod_3426_inner, "mod_3426");
    Operation_IFC mod_3427_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3427 <- mkDebugOperation(mod_3427_inner, "mod_3427");
    Operation_IFC mod_3428_inner <- mkUnaryMap(1713, silu_tile);
    Operation_IFC mod_3428 <- mkDebugOperation(mod_3428_inner, "mod_3428");
    Operation_IFC mod_3429_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3429 <- mkDebugOperation(mod_3429_inner, "mod_3429");
    Operation_IFC mod_3430_inner <- mkBinaryMap(1585, matmul_t_tile);
    Operation_IFC mod_3430 <- mkDebugOperation(mod_3430_inner, "mod_3430");
    PMU_IFC mod_3431_bufferize <- mkPMU(2);
    Operation_IFC mod_3431_inner = mod_3431_bufferize.operation;
    Operation_IFC mod_3431 <- mkDebugOperation(mod_3431_inner, "mod_3431");
    Operation_IFC mod_3432_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3432 <- mkDebugOperation(mod_3432_inner, "mod_3432");
    Operation_IFC mod_3433_inner <- mkFlatten(1);
    Operation_IFC mod_3433 <- mkDebugOperation(mod_3433_inner, "mod_3433");
    Operation_IFC mod_3434_inner <- mkFlatten(0);
    Operation_IFC mod_3434 <- mkDebugOperation(mod_3434_inner, "mod_3434");
    PMU_IFC mod_3435_bufferize <- mkPMU(1);
    Operation_IFC mod_3435_inner = mod_3435_bufferize.operation;
    Operation_IFC mod_3435 <- mkDebugOperation(mod_3435_inner, "mod_3435");
    Operation_IFC mod_3436_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3436 <- mkDebugOperation(mod_3436_inner, "mod_3436");
    PMU_IFC mod_3437_bufferize <- mkPMU(2);
    Operation_IFC mod_3437_inner = mod_3437_bufferize.operation;
    Operation_IFC mod_3437 <- mkDebugOperation(mod_3437_inner, "mod_3437");
    Operation_IFC mod_3438_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3438 <- mkDebugOperation(mod_3438_inner, "mod_3438");
    Operation_IFC mod_3439_inner <- mkFlatten(1);
    Operation_IFC mod_3439 <- mkDebugOperation(mod_3439_inner, "mod_3439");
    Operation_IFC mod_3440_inner <- mkFlatten(0);
    Operation_IFC mod_3440 <- mkDebugOperation(mod_3440_inner, "mod_3440");
    Operation_IFC mod_3441_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3441 <- mkDebugOperation(mod_3441_inner, "mod_3441");
    Operation_IFC mod_3442_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3442 <- mkDebugOperation(mod_3442_inner, "mod_3442");
    PMU_IFC mod_3443_bufferize <- mkPMU(2);
    Operation_IFC mod_3443_inner = mod_3443_bufferize.operation;
    Operation_IFC mod_3443 <- mkDebugOperation(mod_3443_inner, "mod_3443");
    rule rule_4400;
        ChannelMessage t;
        t <- mod_3413.get(0);
        mod_3414.put(0, t);
    endrule
    rule rule_4401;
        ChannelMessage t;
        t <- mod_3409.get(0);
        mod_3442.put(0, t);
    endrule
    rule rule_4402;
        ChannelMessage t;
        t <- mod_3442.get(0);
        mod_3409.put(1, t);
    endrule
    rule rule_4403;
        ChannelMessage t;
        t <- mod_3443.get(1);
        mod_3407.put(1, t);
    endrule
    rule rule_4404;
        ChannelMessage t;
        t <- mod_3412.get(0);
        mod_3413.put(0, t);
    endrule
    rule rule_4405;
        ChannelMessage t;
        t <- mod_3424.get(0);
        mod_3423.put(1, t);
    endrule
    rule rule_4406;
        ChannelMessage t;
        t <- mod_3435.get(0);
        mod_3436.put(0, t);
    endrule
    rule rule_4407;
        ChannelMessage t;
        t <- mod_3435.get(1);
        mod_3430.put(0, t);
    endrule
    rule rule_4408;
        ChannelMessage t;
        t <- mod_3423.get(0);
        mod_3424.put(0, t);
    endrule
    rule rule_4409;
        ChannelMessage t;
        t <- mod_3418.get(0);
        mod_3422.put(0, t);
    endrule
    rule rule_4410;
        ChannelMessage t;
        t <- mod_3418.get(1);
        mod_3419.put(0, t);
    endrule
    rule rule_4411;
        ChannelMessage t;
        t <- mod_3430.get(0);
        mod_3429.put(0, t);
    endrule
    rule rule_4412;
        ChannelMessage t;
        t <- mod_3429.get(0);
        mod_3428.put(0, t);
    endrule
    rule rule_4413;
        ChannelMessage t;
        t <- mod_3437.get(0);
        mod_3438.put(0, t);
    endrule
    rule rule_4414;
        ChannelMessage t;
        t <- mod_3431.get(1);
        mod_3430.put(1, t);
    endrule
    rule rule_4415;
        ChannelMessage t;
        t <- mod_3415.get(1);
        mod_3416.put(0, t);
    endrule
    rule rule_4416;
        ChannelMessage t;
        t <- mod_3410.get(0);
        mod_3435.put(0, t);
    endrule
    rule rule_4417;
        ChannelMessage t;
        t <- mod_3439.get(0);
        mod_3437.put(0, t);
    endrule
    rule rule_4418;
        ChannelMessage t;
        t <- mod_3443.get(0);
        mod_3443.put(1, t);
    endrule
    rule rule_4419;
        ChannelMessage t;
        t <- mod_3414.get(0);
        mod_3415.put(0, t);
    endrule
    rule rule_4420;
        ChannelMessage t;
        t <- mod_3411.get(0);
        mod_3441.put(0, t);
    endrule
    rule rule_4421;
        ChannelMessage t;
        t <- mod_3427.get(0);
        mod_3415.put(1, t);
    endrule
    rule rule_4422;
        ChannelMessage t;
        t <- mod_3433.get(0);
        mod_3431.put(0, t);
    endrule
    rule rule_4423;
        ChannelMessage t;
        t <- mod_3437.get(1);
        mod_3412.put(1, t);
    endrule
    rule rule_4424;
        ChannelMessage t;
        t <- mod_3434.get(0);
        mod_3433.put(0, t);
    endrule
    rule rule_4425;
        ChannelMessage t;
        t <- mod_3440.get(0);
        mod_3439.put(0, t);
    endrule
    rule rule_4426;
        ChannelMessage t;
        t <- mod_3416.get(0);
        mod_3417.put(0, t);
    endrule
    rule rule_4427;
        ChannelMessage t;
        t <- mod_3405.get(0);
        mod_3406.put(0, t);
    endrule
    rule rule_4428;
        ChannelMessage t;
        t <- mod_3423.get(1);
        mod_3416.put(1, t);
    endrule
    rule rule_4429;
        ChannelMessage t;
        t <- mod_3421.get(1);
        mod_3419.put(1, t);
    endrule
    rule rule_4430;
        ChannelMessage t;
        t <- mod_3431.get(0);
        mod_3432.put(0, t);
    endrule
    rule rule_4431;
        ChannelMessage t;
        t <- mod_3410.get(1);
        mod_3411.put(0, t);
    endrule
    rule rule_4432;
        ChannelMessage t;
        t <- mod_3407.get(0);
        mod_3443.put(0, t);
    endrule
    rule rule_4433;
        ChannelMessage t;
        t <- mod_3409.get(1);
        mod_3410.put(0, t);
    endrule
    rule rule_4434;
        ChannelMessage t;
        t <- mod_3432.get(0);
        mod_3431.put(1, t);
    endrule
    rule rule_4435;
        ChannelMessage t;
        t <- mod_3436.get(0);
        mod_3435.put(1, t);
    endrule
    rule rule_4436;
        ChannelMessage t;
        t <- mod_3425.get(0);
        mod_3423.put(0, t);
    endrule
    rule rule_4437;
        ChannelMessage t;
        t <- mod_3411.get(1);
        mod_3412.put(0, t);
    endrule
    rule rule_4438;
        ChannelMessage t;
        t <- mod_3428.get(0);
        mod_3414.put(1, t);
    endrule
    rule rule_4439;
        ChannelMessage t;
        t <- mod_3438.get(0);
        mod_3437.put(1, t);
    endrule
    rule rule_4440;
        ChannelMessage t;
        t <- mod_3404.get(0);
        mod_3405.put(0, t);
    endrule
    rule rule_4441;
        ChannelMessage t;
        t <- mod_3422.get(1);
        mod_3418.put(1, t);
    endrule
    rule rule_4442;
        ChannelMessage t;
        t <- mod_3419.get(0);
        mod_3421.put(0, t);
    endrule
    rule rule_4443;
        ChannelMessage t;
        t <- mod_3408.get(3);
        mod_3409.put(0, t);
    endrule
    rule rule_4444;
        ChannelMessage t;
        t <- mod_3441.get(0);
        mod_3411.put(1, t);
    endrule
    rule rule_4445;
        ChannelMessage t;
        t <- mod_3415.get(0);
        mod_3427.put(0, t);
    endrule
    rule rule_4446;
        ChannelMessage t;
        t <- mod_3407.get(1);
        mod_3408.put(0, t);
    endrule
    rule rule_4447;
        ChannelMessage t;
        t <- mod_3422.get(0);
        mod_3422.put(1, t);
    endrule
    rule rule_4448;
        ChannelMessage t;
        t <- mod_3421.get(0);
        mod_3421.put(1, t);
    endrule
    rule rule_4449;
        ChannelMessage t;
        t <- mod_3426.get(0);
        mod_3425.put(0, t);
    endrule
    rule rule_4450;
        ChannelMessage t;
        t <- mod_3417.get(0);
        mod_3418.put(0, t);
    endrule
    rule rule_4451;
        ChannelMessage t;
        t <- mod_3419.get(1);
        mod_3420.put(1, t);
    endrule
    rule rule_4452;
        ChannelMessage t;
        t <- mod_3406.get(0);
        mod_3407.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3404.put(0, t);
        end
        if (i == 1) begin
            mod_3420.put(0, t);
        end
        if (i == 2) begin
            mod_3426.put(0, t);
        end
        if (i == 3) begin
            mod_3434.put(0, t);
        end
        if (i == 4) begin
            mod_3440.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_3408.get(0);
        end
        if (i == 3) begin
            t <- mod_3408.get(1);
        end
        if (i == 1) begin
            t <- mod_3408.get(2);
        end
        if (i == 2) begin
            t <- mod_3420.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6118 (Operation_IFC);
    Operation_IFC mod_3445_inner <- mkReshape(2, 64);
    Operation_IFC mod_3445 <- mkDebugOperation(mod_3445_inner, "mod_3445");
    Operation_IFC mod_3446_inner <- mkFlatten(1);
    Operation_IFC mod_3446 <- mkDebugOperation(mod_3446_inner, "mod_3446");
    Operation_IFC mod_3447_inner <- mkFlatten(2);
    Operation_IFC mod_3447 <- mkDebugOperation(mod_3447_inner, "mod_3447");
    Operation_IFC mod_3448_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3448 <- mkDebugOperation(mod_3448_inner, "mod_3448");
    Broadcast_IFC#(4) mod_3449_inner <- mkBroadcast(4);
    Operation_IFC mod_3449 <- mkDebugOperation(mod_3449_inner.op, "mod_3449");
    PMU_IFC mod_3450_bufferize <- mkPMU(2);
    Operation_IFC mod_3450_inner = mod_3450_bufferize.operation;
    Operation_IFC mod_3450 <- mkDebugOperation(mod_3450_inner, "mod_3450");
    Broadcast_IFC#(2) mod_3451_inner <- mkBroadcast(2);
    Operation_IFC mod_3451 <- mkDebugOperation(mod_3451_inner.op, "mod_3451");
    PMU_IFC mod_3452_bufferize <- mkPMU(1);
    Operation_IFC mod_3452_inner = mod_3452_bufferize.operation;
    Operation_IFC mod_3452 <- mkDebugOperation(mod_3452_inner, "mod_3452");
    Operation_IFC mod_3453_inner <- mkBinaryMap(1072, matmul_t_tile);
    Operation_IFC mod_3453 <- mkDebugOperation(mod_3453_inner, "mod_3453");
    Operation_IFC mod_3454_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3454 <- mkDebugOperation(mod_3454_inner, "mod_3454");
    Operation_IFC mod_3455_inner <- mkBinaryMap(1840, mul_tile);
    Operation_IFC mod_3455 <- mkDebugOperation(mod_3455_inner, "mod_3455");
    PMU_IFC mod_3456_bufferize <- mkPMU(1);
    Operation_IFC mod_3456_inner = mod_3456_bufferize.operation;
    Operation_IFC mod_3456 <- mkDebugOperation(mod_3456_inner, "mod_3456");
    Operation_IFC mod_3457_inner <- mkBinaryMap(2395, matmul_t_tile);
    Operation_IFC mod_3457 <- mkDebugOperation(mod_3457_inner, "mod_3457");
    Operation_IFC mod_3458_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3458 <- mkDebugOperation(mod_3458_inner, "mod_3458");
    Operation_IFC mod_3459_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3459 <- mkDebugOperation(mod_3459_inner, "mod_3459");
    Operation_IFC mod_3460_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3460 <- mkDebugOperation(mod_3460_inner, "mod_3460");
    Operation_IFC mod_3461_inner <- mkBinaryMap(2739, mul_tile);
    Operation_IFC mod_3461 <- mkDebugOperation(mod_3461_inner, "mod_3461");
    PMU_IFC mod_3462_bufferize <- mkPMU(1);
    Operation_IFC mod_3462_inner = mod_3462_bufferize.operation;
    Operation_IFC mod_3462 <- mkDebugOperation(mod_3462_inner, "mod_3462");
    PMU_IFC mod_3463_bufferize <- mkPMU(2);
    Operation_IFC mod_3463_inner = mod_3463_bufferize.operation;
    Operation_IFC mod_3463 <- mkDebugOperation(mod_3463_inner, "mod_3463");
    PMU_IFC mod_3464_bufferize <- mkPMU(2);
    Operation_IFC mod_3464_inner = mod_3464_bufferize.operation;
    Operation_IFC mod_3464 <- mkDebugOperation(mod_3464_inner, "mod_3464");
    Operation_IFC mod_3465_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3465 <- mkDebugOperation(mod_3465_inner, "mod_3465");
    Operation_IFC mod_3466_inner <- mkFlatten(1);
    Operation_IFC mod_3466 <- mkDebugOperation(mod_3466_inner, "mod_3466");
    Operation_IFC mod_3467_inner <- mkFlatten(0);
    Operation_IFC mod_3467 <- mkDebugOperation(mod_3467_inner, "mod_3467");
    Operation_IFC mod_3468_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3468 <- mkDebugOperation(mod_3468_inner, "mod_3468");
    Operation_IFC mod_3469_inner <- mkUnaryMap(1712, silu_tile);
    Operation_IFC mod_3469 <- mkDebugOperation(mod_3469_inner, "mod_3469");
    Operation_IFC mod_3470_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3470 <- mkDebugOperation(mod_3470_inner, "mod_3470");
    Operation_IFC mod_3471_inner <- mkBinaryMap(1584, matmul_t_tile);
    Operation_IFC mod_3471 <- mkDebugOperation(mod_3471_inner, "mod_3471");
    PMU_IFC mod_3472_bufferize <- mkPMU(2);
    Operation_IFC mod_3472_inner = mod_3472_bufferize.operation;
    Operation_IFC mod_3472 <- mkDebugOperation(mod_3472_inner, "mod_3472");
    Operation_IFC mod_3473_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3473 <- mkDebugOperation(mod_3473_inner, "mod_3473");
    Operation_IFC mod_3474_inner <- mkFlatten(1);
    Operation_IFC mod_3474 <- mkDebugOperation(mod_3474_inner, "mod_3474");
    Operation_IFC mod_3475_inner <- mkFlatten(0);
    Operation_IFC mod_3475 <- mkDebugOperation(mod_3475_inner, "mod_3475");
    PMU_IFC mod_3476_bufferize <- mkPMU(1);
    Operation_IFC mod_3476_inner = mod_3476_bufferize.operation;
    Operation_IFC mod_3476 <- mkDebugOperation(mod_3476_inner, "mod_3476");
    Operation_IFC mod_3477_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3477 <- mkDebugOperation(mod_3477_inner, "mod_3477");
    PMU_IFC mod_3478_bufferize <- mkPMU(2);
    Operation_IFC mod_3478_inner = mod_3478_bufferize.operation;
    Operation_IFC mod_3478 <- mkDebugOperation(mod_3478_inner, "mod_3478");
    Operation_IFC mod_3479_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3479 <- mkDebugOperation(mod_3479_inner, "mod_3479");
    Operation_IFC mod_3480_inner <- mkFlatten(1);
    Operation_IFC mod_3480 <- mkDebugOperation(mod_3480_inner, "mod_3480");
    Operation_IFC mod_3481_inner <- mkFlatten(0);
    Operation_IFC mod_3481 <- mkDebugOperation(mod_3481_inner, "mod_3481");
    Operation_IFC mod_3482_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3482 <- mkDebugOperation(mod_3482_inner, "mod_3482");
    Operation_IFC mod_3483_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3483 <- mkDebugOperation(mod_3483_inner, "mod_3483");
    PMU_IFC mod_3484_bufferize <- mkPMU(2);
    Operation_IFC mod_3484_inner = mod_3484_bufferize.operation;
    Operation_IFC mod_3484 <- mkDebugOperation(mod_3484_inner, "mod_3484");
    rule rule_4453;
        ChannelMessage t;
        t <- mod_3454.get(0);
        mod_3455.put(0, t);
    endrule
    rule rule_4454;
        ChannelMessage t;
        t <- mod_3452.get(1);
        mod_3453.put(0, t);
    endrule
    rule rule_4455;
        ChannelMessage t;
        t <- mod_3458.get(0);
        mod_3459.put(0, t);
    endrule
    rule rule_4456;
        ChannelMessage t;
        t <- mod_3478.get(1);
        mod_3453.put(1, t);
    endrule
    rule rule_4457;
        ChannelMessage t;
        t <- mod_3476.get(1);
        mod_3471.put(0, t);
    endrule
    rule rule_4458;
        ChannelMessage t;
        t <- mod_3463.get(0);
        mod_3463.put(1, t);
    endrule
    rule rule_4459;
        ChannelMessage t;
        t <- mod_3470.get(0);
        mod_3469.put(0, t);
    endrule
    rule rule_4460;
        ChannelMessage t;
        t <- mod_3456.get(1);
        mod_3457.put(0, t);
    endrule
    rule rule_4461;
        ChannelMessage t;
        t <- mod_3453.get(0);
        mod_3454.put(0, t);
    endrule
    rule rule_4462;
        ChannelMessage t;
        t <- mod_3450.get(0);
        mod_3483.put(0, t);
    endrule
    rule rule_4463;
        ChannelMessage t;
        t <- mod_3445.get(0);
        mod_3446.put(0, t);
    endrule
    rule rule_4464;
        ChannelMessage t;
        t <- mod_3449.get(3);
        mod_3450.put(0, t);
    endrule
    rule rule_4465;
        ChannelMessage t;
        t <- mod_3451.get(1);
        mod_3452.put(0, t);
    endrule
    rule rule_4466;
        ChannelMessage t;
        t <- mod_3460.get(0);
        mod_3462.put(0, t);
    endrule
    rule rule_4467;
        ChannelMessage t;
        t <- mod_3460.get(1);
        mod_3461.put(1, t);
    endrule
    rule rule_4468;
        ChannelMessage t;
        t <- mod_3457.get(0);
        mod_3458.put(0, t);
    endrule
    rule rule_4469;
        ChannelMessage t;
        t <- mod_3475.get(0);
        mod_3474.put(0, t);
    endrule
    rule rule_4470;
        ChannelMessage t;
        t <- mod_3484.get(1);
        mod_3448.put(1, t);
    endrule
    rule rule_4471;
        ChannelMessage t;
        t <- mod_3472.get(0);
        mod_3473.put(0, t);
    endrule
    rule rule_4472;
        ChannelMessage t;
        t <- mod_3482.get(0);
        mod_3452.put(1, t);
    endrule
    rule rule_4473;
        ChannelMessage t;
        t <- mod_3459.get(0);
        mod_3463.put(0, t);
    endrule
    rule rule_4474;
        ChannelMessage t;
        t <- mod_3481.get(0);
        mod_3480.put(0, t);
    endrule
    rule rule_4475;
        ChannelMessage t;
        t <- mod_3477.get(0);
        mod_3476.put(1, t);
    endrule
    rule rule_4476;
        ChannelMessage t;
        t <- mod_3466.get(0);
        mod_3464.put(0, t);
    endrule
    rule rule_4477;
        ChannelMessage t;
        t <- mod_3476.get(0);
        mod_3477.put(0, t);
    endrule
    rule rule_4478;
        ChannelMessage t;
        t <- mod_3456.get(0);
        mod_3468.put(0, t);
    endrule
    rule rule_4479;
        ChannelMessage t;
        t <- mod_3459.get(1);
        mod_3460.put(0, t);
    endrule
    rule rule_4480;
        ChannelMessage t;
        t <- mod_3468.get(0);
        mod_3456.put(1, t);
    endrule
    rule rule_4481;
        ChannelMessage t;
        t <- mod_3452.get(0);
        mod_3482.put(0, t);
    endrule
    rule rule_4482;
        ChannelMessage t;
        t <- mod_3462.get(1);
        mod_3460.put(1, t);
    endrule
    rule rule_4483;
        ChannelMessage t;
        t <- mod_3471.get(0);
        mod_3470.put(0, t);
    endrule
    rule rule_4484;
        ChannelMessage t;
        t <- mod_3465.get(0);
        mod_3464.put(1, t);
    endrule
    rule rule_4485;
        ChannelMessage t;
        t <- mod_3455.get(0);
        mod_3456.put(0, t);
    endrule
    rule rule_4486;
        ChannelMessage t;
        t <- mod_3472.get(1);
        mod_3471.put(1, t);
    endrule
    rule rule_4487;
        ChannelMessage t;
        t <- mod_3447.get(0);
        mod_3448.put(0, t);
    endrule
    rule rule_4488;
        ChannelMessage t;
        t <- mod_3469.get(0);
        mod_3455.put(1, t);
    endrule
    rule rule_4489;
        ChannelMessage t;
        t <- mod_3474.get(0);
        mod_3472.put(0, t);
    endrule
    rule rule_4490;
        ChannelMessage t;
        t <- mod_3464.get(1);
        mod_3457.put(1, t);
    endrule
    rule rule_4491;
        ChannelMessage t;
        t <- mod_3451.get(0);
        mod_3476.put(0, t);
    endrule
    rule rule_4492;
        ChannelMessage t;
        t <- mod_3448.get(1);
        mod_3449.put(0, t);
    endrule
    rule rule_4493;
        ChannelMessage t;
        t <- mod_3446.get(0);
        mod_3447.put(0, t);
    endrule
    rule rule_4494;
        ChannelMessage t;
        t <- mod_3467.get(0);
        mod_3466.put(0, t);
    endrule
    rule rule_4495;
        ChannelMessage t;
        t <- mod_3479.get(0);
        mod_3478.put(1, t);
    endrule
    rule rule_4496;
        ChannelMessage t;
        t <- mod_3450.get(1);
        mod_3451.put(0, t);
    endrule
    rule rule_4497;
        ChannelMessage t;
        t <- mod_3448.get(0);
        mod_3484.put(0, t);
    endrule
    rule rule_4498;
        ChannelMessage t;
        t <- mod_3473.get(0);
        mod_3472.put(1, t);
    endrule
    rule rule_4499;
        ChannelMessage t;
        t <- mod_3464.get(0);
        mod_3465.put(0, t);
    endrule
    rule rule_4500;
        ChannelMessage t;
        t <- mod_3480.get(0);
        mod_3478.put(0, t);
    endrule
    rule rule_4501;
        ChannelMessage t;
        t <- mod_3478.get(0);
        mod_3479.put(0, t);
    endrule
    rule rule_4502;
        ChannelMessage t;
        t <- mod_3484.get(0);
        mod_3484.put(1, t);
    endrule
    rule rule_4503;
        ChannelMessage t;
        t <- mod_3463.get(1);
        mod_3459.put(1, t);
    endrule
    rule rule_4504;
        ChannelMessage t;
        t <- mod_3483.get(0);
        mod_3450.put(1, t);
    endrule
    rule rule_4505;
        ChannelMessage t;
        t <- mod_3462.get(0);
        mod_3462.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3445.put(0, t);
        end
        if (i == 1) begin
            mod_3461.put(0, t);
        end
        if (i == 2) begin
            mod_3467.put(0, t);
        end
        if (i == 3) begin
            mod_3475.put(0, t);
        end
        if (i == 4) begin
            mod_3481.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_3449.get(0);
        end
        if (i == 0) begin
            t <- mod_3449.get(1);
        end
        if (i == 3) begin
            t <- mod_3449.get(2);
        end
        if (i == 2) begin
            t <- mod_3461.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6119 (Operation_IFC);
    Operation_IFC mod_3486_inner <- mkReshape(2, 64);
    Operation_IFC mod_3486 <- mkDebugOperation(mod_3486_inner, "mod_3486");
    Operation_IFC mod_3487_inner <- mkFlatten(1);
    Operation_IFC mod_3487 <- mkDebugOperation(mod_3487_inner, "mod_3487");
    Operation_IFC mod_3488_inner <- mkFlatten(2);
    Operation_IFC mod_3488 <- mkDebugOperation(mod_3488_inner, "mod_3488");
    Operation_IFC mod_3489_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3489 <- mkDebugOperation(mod_3489_inner, "mod_3489");
    Broadcast_IFC#(4) mod_3490_inner <- mkBroadcast(4);
    Operation_IFC mod_3490 <- mkDebugOperation(mod_3490_inner.op, "mod_3490");
    PMU_IFC mod_3491_bufferize <- mkPMU(2);
    Operation_IFC mod_3491_inner = mod_3491_bufferize.operation;
    Operation_IFC mod_3491 <- mkDebugOperation(mod_3491_inner, "mod_3491");
    Broadcast_IFC#(2) mod_3492_inner <- mkBroadcast(2);
    Operation_IFC mod_3492 <- mkDebugOperation(mod_3492_inner.op, "mod_3492");
    PMU_IFC mod_3493_bufferize <- mkPMU(1);
    Operation_IFC mod_3493_inner = mod_3493_bufferize.operation;
    Operation_IFC mod_3493 <- mkDebugOperation(mod_3493_inner, "mod_3493");
    Operation_IFC mod_3494_inner <- mkBinaryMap(1071, matmul_t_tile);
    Operation_IFC mod_3494 <- mkDebugOperation(mod_3494_inner, "mod_3494");
    Operation_IFC mod_3495_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3495 <- mkDebugOperation(mod_3495_inner, "mod_3495");
    Operation_IFC mod_3496_inner <- mkBinaryMap(1839, mul_tile);
    Operation_IFC mod_3496 <- mkDebugOperation(mod_3496_inner, "mod_3496");
    PMU_IFC mod_3497_bufferize <- mkPMU(1);
    Operation_IFC mod_3497_inner = mod_3497_bufferize.operation;
    Operation_IFC mod_3497 <- mkDebugOperation(mod_3497_inner, "mod_3497");
    Operation_IFC mod_3498_inner <- mkBinaryMap(2393, matmul_t_tile);
    Operation_IFC mod_3498 <- mkDebugOperation(mod_3498_inner, "mod_3498");
    Operation_IFC mod_3499_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3499 <- mkDebugOperation(mod_3499_inner, "mod_3499");
    Operation_IFC mod_3500_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3500 <- mkDebugOperation(mod_3500_inner, "mod_3500");
    Operation_IFC mod_3501_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3501 <- mkDebugOperation(mod_3501_inner, "mod_3501");
    Operation_IFC mod_3502_inner <- mkBinaryMap(2738, mul_tile);
    Operation_IFC mod_3502 <- mkDebugOperation(mod_3502_inner, "mod_3502");
    PMU_IFC mod_3503_bufferize <- mkPMU(1);
    Operation_IFC mod_3503_inner = mod_3503_bufferize.operation;
    Operation_IFC mod_3503 <- mkDebugOperation(mod_3503_inner, "mod_3503");
    PMU_IFC mod_3504_bufferize <- mkPMU(2);
    Operation_IFC mod_3504_inner = mod_3504_bufferize.operation;
    Operation_IFC mod_3504 <- mkDebugOperation(mod_3504_inner, "mod_3504");
    PMU_IFC mod_3505_bufferize <- mkPMU(2);
    Operation_IFC mod_3505_inner = mod_3505_bufferize.operation;
    Operation_IFC mod_3505 <- mkDebugOperation(mod_3505_inner, "mod_3505");
    Operation_IFC mod_3506_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3506 <- mkDebugOperation(mod_3506_inner, "mod_3506");
    Operation_IFC mod_3507_inner <- mkFlatten(1);
    Operation_IFC mod_3507 <- mkDebugOperation(mod_3507_inner, "mod_3507");
    Operation_IFC mod_3508_inner <- mkFlatten(0);
    Operation_IFC mod_3508 <- mkDebugOperation(mod_3508_inner, "mod_3508");
    Operation_IFC mod_3509_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3509 <- mkDebugOperation(mod_3509_inner, "mod_3509");
    Operation_IFC mod_3510_inner <- mkUnaryMap(1711, silu_tile);
    Operation_IFC mod_3510 <- mkDebugOperation(mod_3510_inner, "mod_3510");
    Operation_IFC mod_3511_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3511 <- mkDebugOperation(mod_3511_inner, "mod_3511");
    Operation_IFC mod_3512_inner <- mkBinaryMap(1583, matmul_t_tile);
    Operation_IFC mod_3512 <- mkDebugOperation(mod_3512_inner, "mod_3512");
    PMU_IFC mod_3513_bufferize <- mkPMU(2);
    Operation_IFC mod_3513_inner = mod_3513_bufferize.operation;
    Operation_IFC mod_3513 <- mkDebugOperation(mod_3513_inner, "mod_3513");
    Operation_IFC mod_3514_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3514 <- mkDebugOperation(mod_3514_inner, "mod_3514");
    Operation_IFC mod_3515_inner <- mkFlatten(1);
    Operation_IFC mod_3515 <- mkDebugOperation(mod_3515_inner, "mod_3515");
    Operation_IFC mod_3516_inner <- mkFlatten(0);
    Operation_IFC mod_3516 <- mkDebugOperation(mod_3516_inner, "mod_3516");
    PMU_IFC mod_3517_bufferize <- mkPMU(1);
    Operation_IFC mod_3517_inner = mod_3517_bufferize.operation;
    Operation_IFC mod_3517 <- mkDebugOperation(mod_3517_inner, "mod_3517");
    Operation_IFC mod_3518_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3518 <- mkDebugOperation(mod_3518_inner, "mod_3518");
    PMU_IFC mod_3519_bufferize <- mkPMU(2);
    Operation_IFC mod_3519_inner = mod_3519_bufferize.operation;
    Operation_IFC mod_3519 <- mkDebugOperation(mod_3519_inner, "mod_3519");
    Operation_IFC mod_3520_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3520 <- mkDebugOperation(mod_3520_inner, "mod_3520");
    Operation_IFC mod_3521_inner <- mkFlatten(1);
    Operation_IFC mod_3521 <- mkDebugOperation(mod_3521_inner, "mod_3521");
    Operation_IFC mod_3522_inner <- mkFlatten(0);
    Operation_IFC mod_3522 <- mkDebugOperation(mod_3522_inner, "mod_3522");
    Operation_IFC mod_3523_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3523 <- mkDebugOperation(mod_3523_inner, "mod_3523");
    Operation_IFC mod_3524_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3524 <- mkDebugOperation(mod_3524_inner, "mod_3524");
    PMU_IFC mod_3525_bufferize <- mkPMU(2);
    Operation_IFC mod_3525_inner = mod_3525_bufferize.operation;
    Operation_IFC mod_3525 <- mkDebugOperation(mod_3525_inner, "mod_3525");
    rule rule_4506;
        ChannelMessage t;
        t <- mod_3492.get(0);
        mod_3517.put(0, t);
    endrule
    rule rule_4507;
        ChannelMessage t;
        t <- mod_3504.get(0);
        mod_3504.put(1, t);
    endrule
    rule rule_4508;
        ChannelMessage t;
        t <- mod_3493.get(1);
        mod_3494.put(0, t);
    endrule
    rule rule_4509;
        ChannelMessage t;
        t <- mod_3517.get(1);
        mod_3512.put(0, t);
    endrule
    rule rule_4510;
        ChannelMessage t;
        t <- mod_3519.get(0);
        mod_3520.put(0, t);
    endrule
    rule rule_4511;
        ChannelMessage t;
        t <- mod_3501.get(1);
        mod_3502.put(1, t);
    endrule
    rule rule_4512;
        ChannelMessage t;
        t <- mod_3514.get(0);
        mod_3513.put(1, t);
    endrule
    rule rule_4513;
        ChannelMessage t;
        t <- mod_3500.get(1);
        mod_3501.put(0, t);
    endrule
    rule rule_4514;
        ChannelMessage t;
        t <- mod_3492.get(1);
        mod_3493.put(0, t);
    endrule
    rule rule_4515;
        ChannelMessage t;
        t <- mod_3491.get(0);
        mod_3524.put(0, t);
    endrule
    rule rule_4516;
        ChannelMessage t;
        t <- mod_3491.get(1);
        mod_3492.put(0, t);
    endrule
    rule rule_4517;
        ChannelMessage t;
        t <- mod_3510.get(0);
        mod_3496.put(1, t);
    endrule
    rule rule_4518;
        ChannelMessage t;
        t <- mod_3495.get(0);
        mod_3496.put(0, t);
    endrule
    rule rule_4519;
        ChannelMessage t;
        t <- mod_3508.get(0);
        mod_3507.put(0, t);
    endrule
    rule rule_4520;
        ChannelMessage t;
        t <- mod_3497.get(0);
        mod_3509.put(0, t);
    endrule
    rule rule_4521;
        ChannelMessage t;
        t <- mod_3519.get(1);
        mod_3494.put(1, t);
    endrule
    rule rule_4522;
        ChannelMessage t;
        t <- mod_3487.get(0);
        mod_3488.put(0, t);
    endrule
    rule rule_4523;
        ChannelMessage t;
        t <- mod_3515.get(0);
        mod_3513.put(0, t);
    endrule
    rule rule_4524;
        ChannelMessage t;
        t <- mod_3490.get(3);
        mod_3491.put(0, t);
    endrule
    rule rule_4525;
        ChannelMessage t;
        t <- mod_3503.get(1);
        mod_3501.put(1, t);
    endrule
    rule rule_4526;
        ChannelMessage t;
        t <- mod_3521.get(0);
        mod_3519.put(0, t);
    endrule
    rule rule_4527;
        ChannelMessage t;
        t <- mod_3524.get(0);
        mod_3491.put(1, t);
    endrule
    rule rule_4528;
        ChannelMessage t;
        t <- mod_3505.get(1);
        mod_3498.put(1, t);
    endrule
    rule rule_4529;
        ChannelMessage t;
        t <- mod_3511.get(0);
        mod_3510.put(0, t);
    endrule
    rule rule_4530;
        ChannelMessage t;
        t <- mod_3494.get(0);
        mod_3495.put(0, t);
    endrule
    rule rule_4531;
        ChannelMessage t;
        t <- mod_3525.get(0);
        mod_3525.put(1, t);
    endrule
    rule rule_4532;
        ChannelMessage t;
        t <- mod_3493.get(0);
        mod_3523.put(0, t);
    endrule
    rule rule_4533;
        ChannelMessage t;
        t <- mod_3509.get(0);
        mod_3497.put(1, t);
    endrule
    rule rule_4534;
        ChannelMessage t;
        t <- mod_3489.get(1);
        mod_3490.put(0, t);
    endrule
    rule rule_4535;
        ChannelMessage t;
        t <- mod_3504.get(1);
        mod_3500.put(1, t);
    endrule
    rule rule_4536;
        ChannelMessage t;
        t <- mod_3525.get(1);
        mod_3489.put(1, t);
    endrule
    rule rule_4537;
        ChannelMessage t;
        t <- mod_3520.get(0);
        mod_3519.put(1, t);
    endrule
    rule rule_4538;
        ChannelMessage t;
        t <- mod_3513.get(1);
        mod_3512.put(1, t);
    endrule
    rule rule_4539;
        ChannelMessage t;
        t <- mod_3497.get(1);
        mod_3498.put(0, t);
    endrule
    rule rule_4540;
        ChannelMessage t;
        t <- mod_3503.get(0);
        mod_3503.put(1, t);
    endrule
    rule rule_4541;
        ChannelMessage t;
        t <- mod_3506.get(0);
        mod_3505.put(1, t);
    endrule
    rule rule_4542;
        ChannelMessage t;
        t <- mod_3517.get(0);
        mod_3518.put(0, t);
    endrule
    rule rule_4543;
        ChannelMessage t;
        t <- mod_3522.get(0);
        mod_3521.put(0, t);
    endrule
    rule rule_4544;
        ChannelMessage t;
        t <- mod_3488.get(0);
        mod_3489.put(0, t);
    endrule
    rule rule_4545;
        ChannelMessage t;
        t <- mod_3500.get(0);
        mod_3504.put(0, t);
    endrule
    rule rule_4546;
        ChannelMessage t;
        t <- mod_3501.get(0);
        mod_3503.put(0, t);
    endrule
    rule rule_4547;
        ChannelMessage t;
        t <- mod_3486.get(0);
        mod_3487.put(0, t);
    endrule
    rule rule_4548;
        ChannelMessage t;
        t <- mod_3516.get(0);
        mod_3515.put(0, t);
    endrule
    rule rule_4549;
        ChannelMessage t;
        t <- mod_3523.get(0);
        mod_3493.put(1, t);
    endrule
    rule rule_4550;
        ChannelMessage t;
        t <- mod_3496.get(0);
        mod_3497.put(0, t);
    endrule
    rule rule_4551;
        ChannelMessage t;
        t <- mod_3507.get(0);
        mod_3505.put(0, t);
    endrule
    rule rule_4552;
        ChannelMessage t;
        t <- mod_3513.get(0);
        mod_3514.put(0, t);
    endrule
    rule rule_4553;
        ChannelMessage t;
        t <- mod_3499.get(0);
        mod_3500.put(0, t);
    endrule
    rule rule_4554;
        ChannelMessage t;
        t <- mod_3512.get(0);
        mod_3511.put(0, t);
    endrule
    rule rule_4555;
        ChannelMessage t;
        t <- mod_3498.get(0);
        mod_3499.put(0, t);
    endrule
    rule rule_4556;
        ChannelMessage t;
        t <- mod_3489.get(0);
        mod_3525.put(0, t);
    endrule
    rule rule_4557;
        ChannelMessage t;
        t <- mod_3505.get(0);
        mod_3506.put(0, t);
    endrule
    rule rule_4558;
        ChannelMessage t;
        t <- mod_3518.get(0);
        mod_3517.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3486.put(0, t);
        end
        if (i == 1) begin
            mod_3502.put(0, t);
        end
        if (i == 2) begin
            mod_3508.put(0, t);
        end
        if (i == 3) begin
            mod_3516.put(0, t);
        end
        if (i == 4) begin
            mod_3522.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_3490.get(0);
        end
        if (i == 2) begin
            t <- mod_3490.get(1);
        end
        if (i == 3) begin
            t <- mod_3490.get(2);
        end
        if (i == 0) begin
            t <- mod_3502.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6120 (Operation_IFC);
    Operation_IFC mod_3527_inner <- mkReshape(2, 64);
    Operation_IFC mod_3527 <- mkDebugOperation(mod_3527_inner, "mod_3527");
    Operation_IFC mod_3528_inner <- mkFlatten(1);
    Operation_IFC mod_3528 <- mkDebugOperation(mod_3528_inner, "mod_3528");
    Operation_IFC mod_3529_inner <- mkFlatten(2);
    Operation_IFC mod_3529 <- mkDebugOperation(mod_3529_inner, "mod_3529");
    Operation_IFC mod_3530_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3530 <- mkDebugOperation(mod_3530_inner, "mod_3530");
    Broadcast_IFC#(4) mod_3531_inner <- mkBroadcast(4);
    Operation_IFC mod_3531 <- mkDebugOperation(mod_3531_inner.op, "mod_3531");
    PMU_IFC mod_3532_bufferize <- mkPMU(2);
    Operation_IFC mod_3532_inner = mod_3532_bufferize.operation;
    Operation_IFC mod_3532 <- mkDebugOperation(mod_3532_inner, "mod_3532");
    Broadcast_IFC#(2) mod_3533_inner <- mkBroadcast(2);
    Operation_IFC mod_3533 <- mkDebugOperation(mod_3533_inner.op, "mod_3533");
    PMU_IFC mod_3534_bufferize <- mkPMU(1);
    Operation_IFC mod_3534_inner = mod_3534_bufferize.operation;
    Operation_IFC mod_3534 <- mkDebugOperation(mod_3534_inner, "mod_3534");
    Operation_IFC mod_3535_inner <- mkBinaryMap(1070, matmul_t_tile);
    Operation_IFC mod_3535 <- mkDebugOperation(mod_3535_inner, "mod_3535");
    Operation_IFC mod_3536_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3536 <- mkDebugOperation(mod_3536_inner, "mod_3536");
    Operation_IFC mod_3537_inner <- mkBinaryMap(1838, mul_tile);
    Operation_IFC mod_3537 <- mkDebugOperation(mod_3537_inner, "mod_3537");
    PMU_IFC mod_3538_bufferize <- mkPMU(1);
    Operation_IFC mod_3538_inner = mod_3538_bufferize.operation;
    Operation_IFC mod_3538 <- mkDebugOperation(mod_3538_inner, "mod_3538");
    Operation_IFC mod_3539_inner <- mkBinaryMap(2391, matmul_t_tile);
    Operation_IFC mod_3539 <- mkDebugOperation(mod_3539_inner, "mod_3539");
    Operation_IFC mod_3540_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3540 <- mkDebugOperation(mod_3540_inner, "mod_3540");
    Operation_IFC mod_3541_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3541 <- mkDebugOperation(mod_3541_inner, "mod_3541");
    Operation_IFC mod_3542_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3542 <- mkDebugOperation(mod_3542_inner, "mod_3542");
    Operation_IFC mod_3543_inner <- mkBinaryMap(2737, mul_tile);
    Operation_IFC mod_3543 <- mkDebugOperation(mod_3543_inner, "mod_3543");
    PMU_IFC mod_3544_bufferize <- mkPMU(1);
    Operation_IFC mod_3544_inner = mod_3544_bufferize.operation;
    Operation_IFC mod_3544 <- mkDebugOperation(mod_3544_inner, "mod_3544");
    PMU_IFC mod_3545_bufferize <- mkPMU(2);
    Operation_IFC mod_3545_inner = mod_3545_bufferize.operation;
    Operation_IFC mod_3545 <- mkDebugOperation(mod_3545_inner, "mod_3545");
    PMU_IFC mod_3546_bufferize <- mkPMU(2);
    Operation_IFC mod_3546_inner = mod_3546_bufferize.operation;
    Operation_IFC mod_3546 <- mkDebugOperation(mod_3546_inner, "mod_3546");
    Operation_IFC mod_3547_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3547 <- mkDebugOperation(mod_3547_inner, "mod_3547");
    Operation_IFC mod_3548_inner <- mkFlatten(1);
    Operation_IFC mod_3548 <- mkDebugOperation(mod_3548_inner, "mod_3548");
    Operation_IFC mod_3549_inner <- mkFlatten(0);
    Operation_IFC mod_3549 <- mkDebugOperation(mod_3549_inner, "mod_3549");
    Operation_IFC mod_3550_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3550 <- mkDebugOperation(mod_3550_inner, "mod_3550");
    Operation_IFC mod_3551_inner <- mkUnaryMap(1710, silu_tile);
    Operation_IFC mod_3551 <- mkDebugOperation(mod_3551_inner, "mod_3551");
    Operation_IFC mod_3552_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3552 <- mkDebugOperation(mod_3552_inner, "mod_3552");
    Operation_IFC mod_3553_inner <- mkBinaryMap(1582, matmul_t_tile);
    Operation_IFC mod_3553 <- mkDebugOperation(mod_3553_inner, "mod_3553");
    PMU_IFC mod_3554_bufferize <- mkPMU(2);
    Operation_IFC mod_3554_inner = mod_3554_bufferize.operation;
    Operation_IFC mod_3554 <- mkDebugOperation(mod_3554_inner, "mod_3554");
    Operation_IFC mod_3555_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3555 <- mkDebugOperation(mod_3555_inner, "mod_3555");
    Operation_IFC mod_3556_inner <- mkFlatten(1);
    Operation_IFC mod_3556 <- mkDebugOperation(mod_3556_inner, "mod_3556");
    Operation_IFC mod_3557_inner <- mkFlatten(0);
    Operation_IFC mod_3557 <- mkDebugOperation(mod_3557_inner, "mod_3557");
    PMU_IFC mod_3558_bufferize <- mkPMU(1);
    Operation_IFC mod_3558_inner = mod_3558_bufferize.operation;
    Operation_IFC mod_3558 <- mkDebugOperation(mod_3558_inner, "mod_3558");
    Operation_IFC mod_3559_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3559 <- mkDebugOperation(mod_3559_inner, "mod_3559");
    PMU_IFC mod_3560_bufferize <- mkPMU(2);
    Operation_IFC mod_3560_inner = mod_3560_bufferize.operation;
    Operation_IFC mod_3560 <- mkDebugOperation(mod_3560_inner, "mod_3560");
    Operation_IFC mod_3561_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3561 <- mkDebugOperation(mod_3561_inner, "mod_3561");
    Operation_IFC mod_3562_inner <- mkFlatten(1);
    Operation_IFC mod_3562 <- mkDebugOperation(mod_3562_inner, "mod_3562");
    Operation_IFC mod_3563_inner <- mkFlatten(0);
    Operation_IFC mod_3563 <- mkDebugOperation(mod_3563_inner, "mod_3563");
    Operation_IFC mod_3564_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3564 <- mkDebugOperation(mod_3564_inner, "mod_3564");
    Operation_IFC mod_3565_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3565 <- mkDebugOperation(mod_3565_inner, "mod_3565");
    PMU_IFC mod_3566_bufferize <- mkPMU(2);
    Operation_IFC mod_3566_inner = mod_3566_bufferize.operation;
    Operation_IFC mod_3566 <- mkDebugOperation(mod_3566_inner, "mod_3566");
    rule rule_4559;
        ChannelMessage t;
        t <- mod_3544.get(0);
        mod_3544.put(1, t);
    endrule
    rule rule_4560;
        ChannelMessage t;
        t <- mod_3530.get(1);
        mod_3531.put(0, t);
    endrule
    rule rule_4561;
        ChannelMessage t;
        t <- mod_3532.get(1);
        mod_3533.put(0, t);
    endrule
    rule rule_4562;
        ChannelMessage t;
        t <- mod_3554.get(0);
        mod_3555.put(0, t);
    endrule
    rule rule_4563;
        ChannelMessage t;
        t <- mod_3554.get(1);
        mod_3553.put(1, t);
    endrule
    rule rule_4564;
        ChannelMessage t;
        t <- mod_3539.get(0);
        mod_3540.put(0, t);
    endrule
    rule rule_4565;
        ChannelMessage t;
        t <- mod_3565.get(0);
        mod_3532.put(1, t);
    endrule
    rule rule_4566;
        ChannelMessage t;
        t <- mod_3563.get(0);
        mod_3562.put(0, t);
    endrule
    rule rule_4567;
        ChannelMessage t;
        t <- mod_3535.get(0);
        mod_3536.put(0, t);
    endrule
    rule rule_4568;
        ChannelMessage t;
        t <- mod_3561.get(0);
        mod_3560.put(1, t);
    endrule
    rule rule_4569;
        ChannelMessage t;
        t <- mod_3549.get(0);
        mod_3548.put(0, t);
    endrule
    rule rule_4570;
        ChannelMessage t;
        t <- mod_3560.get(0);
        mod_3561.put(0, t);
    endrule
    rule rule_4571;
        ChannelMessage t;
        t <- mod_3545.get(1);
        mod_3541.put(1, t);
    endrule
    rule rule_4572;
        ChannelMessage t;
        t <- mod_3562.get(0);
        mod_3560.put(0, t);
    endrule
    rule rule_4573;
        ChannelMessage t;
        t <- mod_3537.get(0);
        mod_3538.put(0, t);
    endrule
    rule rule_4574;
        ChannelMessage t;
        t <- mod_3541.get(0);
        mod_3545.put(0, t);
    endrule
    rule rule_4575;
        ChannelMessage t;
        t <- mod_3542.get(0);
        mod_3544.put(0, t);
    endrule
    rule rule_4576;
        ChannelMessage t;
        t <- mod_3555.get(0);
        mod_3554.put(1, t);
    endrule
    rule rule_4577;
        ChannelMessage t;
        t <- mod_3528.get(0);
        mod_3529.put(0, t);
    endrule
    rule rule_4578;
        ChannelMessage t;
        t <- mod_3559.get(0);
        mod_3558.put(1, t);
    endrule
    rule rule_4579;
        ChannelMessage t;
        t <- mod_3552.get(0);
        mod_3551.put(0, t);
    endrule
    rule rule_4580;
        ChannelMessage t;
        t <- mod_3544.get(1);
        mod_3542.put(1, t);
    endrule
    rule rule_4581;
        ChannelMessage t;
        t <- mod_3534.get(1);
        mod_3535.put(0, t);
    endrule
    rule rule_4582;
        ChannelMessage t;
        t <- mod_3530.get(0);
        mod_3566.put(0, t);
    endrule
    rule rule_4583;
        ChannelMessage t;
        t <- mod_3550.get(0);
        mod_3538.put(1, t);
    endrule
    rule rule_4584;
        ChannelMessage t;
        t <- mod_3553.get(0);
        mod_3552.put(0, t);
    endrule
    rule rule_4585;
        ChannelMessage t;
        t <- mod_3566.get(1);
        mod_3530.put(1, t);
    endrule
    rule rule_4586;
        ChannelMessage t;
        t <- mod_3533.get(0);
        mod_3558.put(0, t);
    endrule
    rule rule_4587;
        ChannelMessage t;
        t <- mod_3540.get(0);
        mod_3541.put(0, t);
    endrule
    rule rule_4588;
        ChannelMessage t;
        t <- mod_3538.get(1);
        mod_3539.put(0, t);
    endrule
    rule rule_4589;
        ChannelMessage t;
        t <- mod_3541.get(1);
        mod_3542.put(0, t);
    endrule
    rule rule_4590;
        ChannelMessage t;
        t <- mod_3546.get(0);
        mod_3547.put(0, t);
    endrule
    rule rule_4591;
        ChannelMessage t;
        t <- mod_3560.get(1);
        mod_3535.put(1, t);
    endrule
    rule rule_4592;
        ChannelMessage t;
        t <- mod_3533.get(1);
        mod_3534.put(0, t);
    endrule
    rule rule_4593;
        ChannelMessage t;
        t <- mod_3564.get(0);
        mod_3534.put(1, t);
    endrule
    rule rule_4594;
        ChannelMessage t;
        t <- mod_3532.get(0);
        mod_3565.put(0, t);
    endrule
    rule rule_4595;
        ChannelMessage t;
        t <- mod_3551.get(0);
        mod_3537.put(1, t);
    endrule
    rule rule_4596;
        ChannelMessage t;
        t <- mod_3566.get(0);
        mod_3566.put(1, t);
    endrule
    rule rule_4597;
        ChannelMessage t;
        t <- mod_3546.get(1);
        mod_3539.put(1, t);
    endrule
    rule rule_4598;
        ChannelMessage t;
        t <- mod_3527.get(0);
        mod_3528.put(0, t);
    endrule
    rule rule_4599;
        ChannelMessage t;
        t <- mod_3534.get(0);
        mod_3564.put(0, t);
    endrule
    rule rule_4600;
        ChannelMessage t;
        t <- mod_3538.get(0);
        mod_3550.put(0, t);
    endrule
    rule rule_4601;
        ChannelMessage t;
        t <- mod_3548.get(0);
        mod_3546.put(0, t);
    endrule
    rule rule_4602;
        ChannelMessage t;
        t <- mod_3557.get(0);
        mod_3556.put(0, t);
    endrule
    rule rule_4603;
        ChannelMessage t;
        t <- mod_3558.get(1);
        mod_3553.put(0, t);
    endrule
    rule rule_4604;
        ChannelMessage t;
        t <- mod_3547.get(0);
        mod_3546.put(1, t);
    endrule
    rule rule_4605;
        ChannelMessage t;
        t <- mod_3558.get(0);
        mod_3559.put(0, t);
    endrule
    rule rule_4606;
        ChannelMessage t;
        t <- mod_3542.get(1);
        mod_3543.put(1, t);
    endrule
    rule rule_4607;
        ChannelMessage t;
        t <- mod_3545.get(0);
        mod_3545.put(1, t);
    endrule
    rule rule_4608;
        ChannelMessage t;
        t <- mod_3529.get(0);
        mod_3530.put(0, t);
    endrule
    rule rule_4609;
        ChannelMessage t;
        t <- mod_3531.get(3);
        mod_3532.put(0, t);
    endrule
    rule rule_4610;
        ChannelMessage t;
        t <- mod_3536.get(0);
        mod_3537.put(0, t);
    endrule
    rule rule_4611;
        ChannelMessage t;
        t <- mod_3556.get(0);
        mod_3554.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3527.put(0, t);
        end
        if (i == 1) begin
            mod_3543.put(0, t);
        end
        if (i == 2) begin
            mod_3549.put(0, t);
        end
        if (i == 3) begin
            mod_3557.put(0, t);
        end
        if (i == 4) begin
            mod_3563.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 2) begin
            t <- mod_3531.get(0);
        end
        if (i == 1) begin
            t <- mod_3531.get(1);
        end
        if (i == 3) begin
            t <- mod_3531.get(2);
        end
        if (i == 0) begin
            t <- mod_3543.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6121 (Operation_IFC);
    Operation_IFC mod_3568_inner <- mkReshape(2, 64);
    Operation_IFC mod_3568 <- mkDebugOperation(mod_3568_inner, "mod_3568");
    Operation_IFC mod_3569_inner <- mkFlatten(1);
    Operation_IFC mod_3569 <- mkDebugOperation(mod_3569_inner, "mod_3569");
    Operation_IFC mod_3570_inner <- mkFlatten(2);
    Operation_IFC mod_3570 <- mkDebugOperation(mod_3570_inner, "mod_3570");
    Operation_IFC mod_3571_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3571 <- mkDebugOperation(mod_3571_inner, "mod_3571");
    Broadcast_IFC#(4) mod_3572_inner <- mkBroadcast(4);
    Operation_IFC mod_3572 <- mkDebugOperation(mod_3572_inner.op, "mod_3572");
    PMU_IFC mod_3573_bufferize <- mkPMU(2);
    Operation_IFC mod_3573_inner = mod_3573_bufferize.operation;
    Operation_IFC mod_3573 <- mkDebugOperation(mod_3573_inner, "mod_3573");
    Broadcast_IFC#(2) mod_3574_inner <- mkBroadcast(2);
    Operation_IFC mod_3574 <- mkDebugOperation(mod_3574_inner.op, "mod_3574");
    PMU_IFC mod_3575_bufferize <- mkPMU(1);
    Operation_IFC mod_3575_inner = mod_3575_bufferize.operation;
    Operation_IFC mod_3575 <- mkDebugOperation(mod_3575_inner, "mod_3575");
    Operation_IFC mod_3576_inner <- mkBinaryMap(1069, matmul_t_tile);
    Operation_IFC mod_3576 <- mkDebugOperation(mod_3576_inner, "mod_3576");
    Operation_IFC mod_3577_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3577 <- mkDebugOperation(mod_3577_inner, "mod_3577");
    Operation_IFC mod_3578_inner <- mkBinaryMap(1837, mul_tile);
    Operation_IFC mod_3578 <- mkDebugOperation(mod_3578_inner, "mod_3578");
    PMU_IFC mod_3579_bufferize <- mkPMU(1);
    Operation_IFC mod_3579_inner = mod_3579_bufferize.operation;
    Operation_IFC mod_3579 <- mkDebugOperation(mod_3579_inner, "mod_3579");
    Operation_IFC mod_3580_inner <- mkBinaryMap(2389, matmul_t_tile);
    Operation_IFC mod_3580 <- mkDebugOperation(mod_3580_inner, "mod_3580");
    Operation_IFC mod_3581_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3581 <- mkDebugOperation(mod_3581_inner, "mod_3581");
    Operation_IFC mod_3582_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3582 <- mkDebugOperation(mod_3582_inner, "mod_3582");
    Operation_IFC mod_3583_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3583 <- mkDebugOperation(mod_3583_inner, "mod_3583");
    Operation_IFC mod_3584_inner <- mkBinaryMap(2736, mul_tile);
    Operation_IFC mod_3584 <- mkDebugOperation(mod_3584_inner, "mod_3584");
    PMU_IFC mod_3585_bufferize <- mkPMU(1);
    Operation_IFC mod_3585_inner = mod_3585_bufferize.operation;
    Operation_IFC mod_3585 <- mkDebugOperation(mod_3585_inner, "mod_3585");
    PMU_IFC mod_3586_bufferize <- mkPMU(2);
    Operation_IFC mod_3586_inner = mod_3586_bufferize.operation;
    Operation_IFC mod_3586 <- mkDebugOperation(mod_3586_inner, "mod_3586");
    PMU_IFC mod_3587_bufferize <- mkPMU(2);
    Operation_IFC mod_3587_inner = mod_3587_bufferize.operation;
    Operation_IFC mod_3587 <- mkDebugOperation(mod_3587_inner, "mod_3587");
    Operation_IFC mod_3588_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3588 <- mkDebugOperation(mod_3588_inner, "mod_3588");
    Operation_IFC mod_3589_inner <- mkFlatten(1);
    Operation_IFC mod_3589 <- mkDebugOperation(mod_3589_inner, "mod_3589");
    Operation_IFC mod_3590_inner <- mkFlatten(0);
    Operation_IFC mod_3590 <- mkDebugOperation(mod_3590_inner, "mod_3590");
    Operation_IFC mod_3591_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3591 <- mkDebugOperation(mod_3591_inner, "mod_3591");
    Operation_IFC mod_3592_inner <- mkUnaryMap(1709, silu_tile);
    Operation_IFC mod_3592 <- mkDebugOperation(mod_3592_inner, "mod_3592");
    Operation_IFC mod_3593_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3593 <- mkDebugOperation(mod_3593_inner, "mod_3593");
    Operation_IFC mod_3594_inner <- mkBinaryMap(1581, matmul_t_tile);
    Operation_IFC mod_3594 <- mkDebugOperation(mod_3594_inner, "mod_3594");
    PMU_IFC mod_3595_bufferize <- mkPMU(2);
    Operation_IFC mod_3595_inner = mod_3595_bufferize.operation;
    Operation_IFC mod_3595 <- mkDebugOperation(mod_3595_inner, "mod_3595");
    Operation_IFC mod_3596_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3596 <- mkDebugOperation(mod_3596_inner, "mod_3596");
    Operation_IFC mod_3597_inner <- mkFlatten(1);
    Operation_IFC mod_3597 <- mkDebugOperation(mod_3597_inner, "mod_3597");
    Operation_IFC mod_3598_inner <- mkFlatten(0);
    Operation_IFC mod_3598 <- mkDebugOperation(mod_3598_inner, "mod_3598");
    PMU_IFC mod_3599_bufferize <- mkPMU(1);
    Operation_IFC mod_3599_inner = mod_3599_bufferize.operation;
    Operation_IFC mod_3599 <- mkDebugOperation(mod_3599_inner, "mod_3599");
    Operation_IFC mod_3600_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3600 <- mkDebugOperation(mod_3600_inner, "mod_3600");
    PMU_IFC mod_3601_bufferize <- mkPMU(2);
    Operation_IFC mod_3601_inner = mod_3601_bufferize.operation;
    Operation_IFC mod_3601 <- mkDebugOperation(mod_3601_inner, "mod_3601");
    Operation_IFC mod_3602_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3602 <- mkDebugOperation(mod_3602_inner, "mod_3602");
    Operation_IFC mod_3603_inner <- mkFlatten(1);
    Operation_IFC mod_3603 <- mkDebugOperation(mod_3603_inner, "mod_3603");
    Operation_IFC mod_3604_inner <- mkFlatten(0);
    Operation_IFC mod_3604 <- mkDebugOperation(mod_3604_inner, "mod_3604");
    Operation_IFC mod_3605_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3605 <- mkDebugOperation(mod_3605_inner, "mod_3605");
    Operation_IFC mod_3606_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3606 <- mkDebugOperation(mod_3606_inner, "mod_3606");
    PMU_IFC mod_3607_bufferize <- mkPMU(2);
    Operation_IFC mod_3607_inner = mod_3607_bufferize.operation;
    Operation_IFC mod_3607 <- mkDebugOperation(mod_3607_inner, "mod_3607");
    rule rule_4612;
        ChannelMessage t;
        t <- mod_3573.get(0);
        mod_3606.put(0, t);
    endrule
    rule rule_4613;
        ChannelMessage t;
        t <- mod_3578.get(0);
        mod_3579.put(0, t);
    endrule
    rule rule_4614;
        ChannelMessage t;
        t <- mod_3598.get(0);
        mod_3597.put(0, t);
    endrule
    rule rule_4615;
        ChannelMessage t;
        t <- mod_3601.get(0);
        mod_3602.put(0, t);
    endrule
    rule rule_4616;
        ChannelMessage t;
        t <- mod_3588.get(0);
        mod_3587.put(1, t);
    endrule
    rule rule_4617;
        ChannelMessage t;
        t <- mod_3571.get(0);
        mod_3607.put(0, t);
    endrule
    rule rule_4618;
        ChannelMessage t;
        t <- mod_3585.get(1);
        mod_3583.put(1, t);
    endrule
    rule rule_4619;
        ChannelMessage t;
        t <- mod_3604.get(0);
        mod_3603.put(0, t);
    endrule
    rule rule_4620;
        ChannelMessage t;
        t <- mod_3586.get(0);
        mod_3586.put(1, t);
    endrule
    rule rule_4621;
        ChannelMessage t;
        t <- mod_3593.get(0);
        mod_3592.put(0, t);
    endrule
    rule rule_4622;
        ChannelMessage t;
        t <- mod_3583.get(0);
        mod_3585.put(0, t);
    endrule
    rule rule_4623;
        ChannelMessage t;
        t <- mod_3587.get(1);
        mod_3580.put(1, t);
    endrule
    rule rule_4624;
        ChannelMessage t;
        t <- mod_3575.get(1);
        mod_3576.put(0, t);
    endrule
    rule rule_4625;
        ChannelMessage t;
        t <- mod_3587.get(0);
        mod_3588.put(0, t);
    endrule
    rule rule_4626;
        ChannelMessage t;
        t <- mod_3589.get(0);
        mod_3587.put(0, t);
    endrule
    rule rule_4627;
        ChannelMessage t;
        t <- mod_3600.get(0);
        mod_3599.put(1, t);
    endrule
    rule rule_4628;
        ChannelMessage t;
        t <- mod_3595.get(0);
        mod_3596.put(0, t);
    endrule
    rule rule_4629;
        ChannelMessage t;
        t <- mod_3573.get(1);
        mod_3574.put(0, t);
    endrule
    rule rule_4630;
        ChannelMessage t;
        t <- mod_3574.get(1);
        mod_3575.put(0, t);
    endrule
    rule rule_4631;
        ChannelMessage t;
        t <- mod_3570.get(0);
        mod_3571.put(0, t);
    endrule
    rule rule_4632;
        ChannelMessage t;
        t <- mod_3579.get(0);
        mod_3591.put(0, t);
    endrule
    rule rule_4633;
        ChannelMessage t;
        t <- mod_3583.get(1);
        mod_3584.put(1, t);
    endrule
    rule rule_4634;
        ChannelMessage t;
        t <- mod_3591.get(0);
        mod_3579.put(1, t);
    endrule
    rule rule_4635;
        ChannelMessage t;
        t <- mod_3575.get(0);
        mod_3605.put(0, t);
    endrule
    rule rule_4636;
        ChannelMessage t;
        t <- mod_3581.get(0);
        mod_3582.put(0, t);
    endrule
    rule rule_4637;
        ChannelMessage t;
        t <- mod_3580.get(0);
        mod_3581.put(0, t);
    endrule
    rule rule_4638;
        ChannelMessage t;
        t <- mod_3605.get(0);
        mod_3575.put(1, t);
    endrule
    rule rule_4639;
        ChannelMessage t;
        t <- mod_3585.get(0);
        mod_3585.put(1, t);
    endrule
    rule rule_4640;
        ChannelMessage t;
        t <- mod_3572.get(3);
        mod_3573.put(0, t);
    endrule
    rule rule_4641;
        ChannelMessage t;
        t <- mod_3597.get(0);
        mod_3595.put(0, t);
    endrule
    rule rule_4642;
        ChannelMessage t;
        t <- mod_3601.get(1);
        mod_3576.put(1, t);
    endrule
    rule rule_4643;
        ChannelMessage t;
        t <- mod_3576.get(0);
        mod_3577.put(0, t);
    endrule
    rule rule_4644;
        ChannelMessage t;
        t <- mod_3596.get(0);
        mod_3595.put(1, t);
    endrule
    rule rule_4645;
        ChannelMessage t;
        t <- mod_3579.get(1);
        mod_3580.put(0, t);
    endrule
    rule rule_4646;
        ChannelMessage t;
        t <- mod_3607.get(1);
        mod_3571.put(1, t);
    endrule
    rule rule_4647;
        ChannelMessage t;
        t <- mod_3599.get(1);
        mod_3594.put(0, t);
    endrule
    rule rule_4648;
        ChannelMessage t;
        t <- mod_3569.get(0);
        mod_3570.put(0, t);
    endrule
    rule rule_4649;
        ChannelMessage t;
        t <- mod_3590.get(0);
        mod_3589.put(0, t);
    endrule
    rule rule_4650;
        ChannelMessage t;
        t <- mod_3592.get(0);
        mod_3578.put(1, t);
    endrule
    rule rule_4651;
        ChannelMessage t;
        t <- mod_3586.get(1);
        mod_3582.put(1, t);
    endrule
    rule rule_4652;
        ChannelMessage t;
        t <- mod_3602.get(0);
        mod_3601.put(1, t);
    endrule
    rule rule_4653;
        ChannelMessage t;
        t <- mod_3568.get(0);
        mod_3569.put(0, t);
    endrule
    rule rule_4654;
        ChannelMessage t;
        t <- mod_3577.get(0);
        mod_3578.put(0, t);
    endrule
    rule rule_4655;
        ChannelMessage t;
        t <- mod_3595.get(1);
        mod_3594.put(1, t);
    endrule
    rule rule_4656;
        ChannelMessage t;
        t <- mod_3571.get(1);
        mod_3572.put(0, t);
    endrule
    rule rule_4657;
        ChannelMessage t;
        t <- mod_3574.get(0);
        mod_3599.put(0, t);
    endrule
    rule rule_4658;
        ChannelMessage t;
        t <- mod_3582.get(0);
        mod_3586.put(0, t);
    endrule
    rule rule_4659;
        ChannelMessage t;
        t <- mod_3607.get(0);
        mod_3607.put(1, t);
    endrule
    rule rule_4660;
        ChannelMessage t;
        t <- mod_3582.get(1);
        mod_3583.put(0, t);
    endrule
    rule rule_4661;
        ChannelMessage t;
        t <- mod_3594.get(0);
        mod_3593.put(0, t);
    endrule
    rule rule_4662;
        ChannelMessage t;
        t <- mod_3599.get(0);
        mod_3600.put(0, t);
    endrule
    rule rule_4663;
        ChannelMessage t;
        t <- mod_3606.get(0);
        mod_3573.put(1, t);
    endrule
    rule rule_4664;
        ChannelMessage t;
        t <- mod_3603.get(0);
        mod_3601.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3568.put(0, t);
        end
        if (i == 1) begin
            mod_3584.put(0, t);
        end
        if (i == 2) begin
            mod_3590.put(0, t);
        end
        if (i == 3) begin
            mod_3598.put(0, t);
        end
        if (i == 4) begin
            mod_3604.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_3572.get(0);
        end
        if (i == 2) begin
            t <- mod_3572.get(1);
        end
        if (i == 3) begin
            t <- mod_3572.get(2);
        end
        if (i == 0) begin
            t <- mod_3584.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6122 (Operation_IFC);
    Operation_IFC mod_3609_inner <- mkReshape(2, 64);
    Operation_IFC mod_3609 <- mkDebugOperation(mod_3609_inner, "mod_3609");
    Operation_IFC mod_3610_inner <- mkFlatten(1);
    Operation_IFC mod_3610 <- mkDebugOperation(mod_3610_inner, "mod_3610");
    Operation_IFC mod_3611_inner <- mkFlatten(2);
    Operation_IFC mod_3611 <- mkDebugOperation(mod_3611_inner, "mod_3611");
    Operation_IFC mod_3612_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3612 <- mkDebugOperation(mod_3612_inner, "mod_3612");
    Broadcast_IFC#(4) mod_3613_inner <- mkBroadcast(4);
    Operation_IFC mod_3613 <- mkDebugOperation(mod_3613_inner.op, "mod_3613");
    PMU_IFC mod_3614_bufferize <- mkPMU(2);
    Operation_IFC mod_3614_inner = mod_3614_bufferize.operation;
    Operation_IFC mod_3614 <- mkDebugOperation(mod_3614_inner, "mod_3614");
    Broadcast_IFC#(2) mod_3615_inner <- mkBroadcast(2);
    Operation_IFC mod_3615 <- mkDebugOperation(mod_3615_inner.op, "mod_3615");
    PMU_IFC mod_3616_bufferize <- mkPMU(1);
    Operation_IFC mod_3616_inner = mod_3616_bufferize.operation;
    Operation_IFC mod_3616 <- mkDebugOperation(mod_3616_inner, "mod_3616");
    Operation_IFC mod_3617_inner <- mkBinaryMap(1068, matmul_t_tile);
    Operation_IFC mod_3617 <- mkDebugOperation(mod_3617_inner, "mod_3617");
    Operation_IFC mod_3618_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3618 <- mkDebugOperation(mod_3618_inner, "mod_3618");
    Operation_IFC mod_3619_inner <- mkBinaryMap(1836, mul_tile);
    Operation_IFC mod_3619 <- mkDebugOperation(mod_3619_inner, "mod_3619");
    PMU_IFC mod_3620_bufferize <- mkPMU(1);
    Operation_IFC mod_3620_inner = mod_3620_bufferize.operation;
    Operation_IFC mod_3620 <- mkDebugOperation(mod_3620_inner, "mod_3620");
    Operation_IFC mod_3621_inner <- mkBinaryMap(2387, matmul_t_tile);
    Operation_IFC mod_3621 <- mkDebugOperation(mod_3621_inner, "mod_3621");
    Operation_IFC mod_3622_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3622 <- mkDebugOperation(mod_3622_inner, "mod_3622");
    Operation_IFC mod_3623_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3623 <- mkDebugOperation(mod_3623_inner, "mod_3623");
    Operation_IFC mod_3624_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3624 <- mkDebugOperation(mod_3624_inner, "mod_3624");
    Operation_IFC mod_3625_inner <- mkBinaryMap(2735, mul_tile);
    Operation_IFC mod_3625 <- mkDebugOperation(mod_3625_inner, "mod_3625");
    PMU_IFC mod_3626_bufferize <- mkPMU(1);
    Operation_IFC mod_3626_inner = mod_3626_bufferize.operation;
    Operation_IFC mod_3626 <- mkDebugOperation(mod_3626_inner, "mod_3626");
    PMU_IFC mod_3627_bufferize <- mkPMU(2);
    Operation_IFC mod_3627_inner = mod_3627_bufferize.operation;
    Operation_IFC mod_3627 <- mkDebugOperation(mod_3627_inner, "mod_3627");
    PMU_IFC mod_3628_bufferize <- mkPMU(2);
    Operation_IFC mod_3628_inner = mod_3628_bufferize.operation;
    Operation_IFC mod_3628 <- mkDebugOperation(mod_3628_inner, "mod_3628");
    Operation_IFC mod_3629_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3629 <- mkDebugOperation(mod_3629_inner, "mod_3629");
    Operation_IFC mod_3630_inner <- mkFlatten(1);
    Operation_IFC mod_3630 <- mkDebugOperation(mod_3630_inner, "mod_3630");
    Operation_IFC mod_3631_inner <- mkFlatten(0);
    Operation_IFC mod_3631 <- mkDebugOperation(mod_3631_inner, "mod_3631");
    Operation_IFC mod_3632_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3632 <- mkDebugOperation(mod_3632_inner, "mod_3632");
    Operation_IFC mod_3633_inner <- mkUnaryMap(1708, silu_tile);
    Operation_IFC mod_3633 <- mkDebugOperation(mod_3633_inner, "mod_3633");
    Operation_IFC mod_3634_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3634 <- mkDebugOperation(mod_3634_inner, "mod_3634");
    Operation_IFC mod_3635_inner <- mkBinaryMap(1580, matmul_t_tile);
    Operation_IFC mod_3635 <- mkDebugOperation(mod_3635_inner, "mod_3635");
    PMU_IFC mod_3636_bufferize <- mkPMU(2);
    Operation_IFC mod_3636_inner = mod_3636_bufferize.operation;
    Operation_IFC mod_3636 <- mkDebugOperation(mod_3636_inner, "mod_3636");
    Operation_IFC mod_3637_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3637 <- mkDebugOperation(mod_3637_inner, "mod_3637");
    Operation_IFC mod_3638_inner <- mkFlatten(1);
    Operation_IFC mod_3638 <- mkDebugOperation(mod_3638_inner, "mod_3638");
    Operation_IFC mod_3639_inner <- mkFlatten(0);
    Operation_IFC mod_3639 <- mkDebugOperation(mod_3639_inner, "mod_3639");
    PMU_IFC mod_3640_bufferize <- mkPMU(1);
    Operation_IFC mod_3640_inner = mod_3640_bufferize.operation;
    Operation_IFC mod_3640 <- mkDebugOperation(mod_3640_inner, "mod_3640");
    Operation_IFC mod_3641_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3641 <- mkDebugOperation(mod_3641_inner, "mod_3641");
    PMU_IFC mod_3642_bufferize <- mkPMU(2);
    Operation_IFC mod_3642_inner = mod_3642_bufferize.operation;
    Operation_IFC mod_3642 <- mkDebugOperation(mod_3642_inner, "mod_3642");
    Operation_IFC mod_3643_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3643 <- mkDebugOperation(mod_3643_inner, "mod_3643");
    Operation_IFC mod_3644_inner <- mkFlatten(1);
    Operation_IFC mod_3644 <- mkDebugOperation(mod_3644_inner, "mod_3644");
    Operation_IFC mod_3645_inner <- mkFlatten(0);
    Operation_IFC mod_3645 <- mkDebugOperation(mod_3645_inner, "mod_3645");
    Operation_IFC mod_3646_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3646 <- mkDebugOperation(mod_3646_inner, "mod_3646");
    Operation_IFC mod_3647_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3647 <- mkDebugOperation(mod_3647_inner, "mod_3647");
    PMU_IFC mod_3648_bufferize <- mkPMU(2);
    Operation_IFC mod_3648_inner = mod_3648_bufferize.operation;
    Operation_IFC mod_3648 <- mkDebugOperation(mod_3648_inner, "mod_3648");
    rule rule_4665;
        ChannelMessage t;
        t <- mod_3620.get(0);
        mod_3632.put(0, t);
    endrule
    rule rule_4666;
        ChannelMessage t;
        t <- mod_3621.get(0);
        mod_3622.put(0, t);
    endrule
    rule rule_4667;
        ChannelMessage t;
        t <- mod_3618.get(0);
        mod_3619.put(0, t);
    endrule
    rule rule_4668;
        ChannelMessage t;
        t <- mod_3624.get(1);
        mod_3625.put(1, t);
    endrule
    rule rule_4669;
        ChannelMessage t;
        t <- mod_3644.get(0);
        mod_3642.put(0, t);
    endrule
    rule rule_4670;
        ChannelMessage t;
        t <- mod_3616.get(0);
        mod_3646.put(0, t);
    endrule
    rule rule_4671;
        ChannelMessage t;
        t <- mod_3642.get(0);
        mod_3643.put(0, t);
    endrule
    rule rule_4672;
        ChannelMessage t;
        t <- mod_3632.get(0);
        mod_3620.put(1, t);
    endrule
    rule rule_4673;
        ChannelMessage t;
        t <- mod_3643.get(0);
        mod_3642.put(1, t);
    endrule
    rule rule_4674;
        ChannelMessage t;
        t <- mod_3629.get(0);
        mod_3628.put(1, t);
    endrule
    rule rule_4675;
        ChannelMessage t;
        t <- mod_3639.get(0);
        mod_3638.put(0, t);
    endrule
    rule rule_4676;
        ChannelMessage t;
        t <- mod_3628.get(0);
        mod_3629.put(0, t);
    endrule
    rule rule_4677;
        ChannelMessage t;
        t <- mod_3614.get(0);
        mod_3647.put(0, t);
    endrule
    rule rule_4678;
        ChannelMessage t;
        t <- mod_3620.get(1);
        mod_3621.put(0, t);
    endrule
    rule rule_4679;
        ChannelMessage t;
        t <- mod_3624.get(0);
        mod_3626.put(0, t);
    endrule
    rule rule_4680;
        ChannelMessage t;
        t <- mod_3613.get(3);
        mod_3614.put(0, t);
    endrule
    rule rule_4681;
        ChannelMessage t;
        t <- mod_3615.get(1);
        mod_3616.put(0, t);
    endrule
    rule rule_4682;
        ChannelMessage t;
        t <- mod_3634.get(0);
        mod_3633.put(0, t);
    endrule
    rule rule_4683;
        ChannelMessage t;
        t <- mod_3645.get(0);
        mod_3644.put(0, t);
    endrule
    rule rule_4684;
        ChannelMessage t;
        t <- mod_3640.get(1);
        mod_3635.put(0, t);
    endrule
    rule rule_4685;
        ChannelMessage t;
        t <- mod_3648.get(1);
        mod_3612.put(1, t);
    endrule
    rule rule_4686;
        ChannelMessage t;
        t <- mod_3609.get(0);
        mod_3610.put(0, t);
    endrule
    rule rule_4687;
        ChannelMessage t;
        t <- mod_3623.get(1);
        mod_3624.put(0, t);
    endrule
    rule rule_4688;
        ChannelMessage t;
        t <- mod_3616.get(1);
        mod_3617.put(0, t);
    endrule
    rule rule_4689;
        ChannelMessage t;
        t <- mod_3626.get(1);
        mod_3624.put(1, t);
    endrule
    rule rule_4690;
        ChannelMessage t;
        t <- mod_3637.get(0);
        mod_3636.put(1, t);
    endrule
    rule rule_4691;
        ChannelMessage t;
        t <- mod_3631.get(0);
        mod_3630.put(0, t);
    endrule
    rule rule_4692;
        ChannelMessage t;
        t <- mod_3647.get(0);
        mod_3614.put(1, t);
    endrule
    rule rule_4693;
        ChannelMessage t;
        t <- mod_3635.get(0);
        mod_3634.put(0, t);
    endrule
    rule rule_4694;
        ChannelMessage t;
        t <- mod_3638.get(0);
        mod_3636.put(0, t);
    endrule
    rule rule_4695;
        ChannelMessage t;
        t <- mod_3619.get(0);
        mod_3620.put(0, t);
    endrule
    rule rule_4696;
        ChannelMessage t;
        t <- mod_3627.get(1);
        mod_3623.put(1, t);
    endrule
    rule rule_4697;
        ChannelMessage t;
        t <- mod_3617.get(0);
        mod_3618.put(0, t);
    endrule
    rule rule_4698;
        ChannelMessage t;
        t <- mod_3646.get(0);
        mod_3616.put(1, t);
    endrule
    rule rule_4699;
        ChannelMessage t;
        t <- mod_3633.get(0);
        mod_3619.put(1, t);
    endrule
    rule rule_4700;
        ChannelMessage t;
        t <- mod_3640.get(0);
        mod_3641.put(0, t);
    endrule
    rule rule_4701;
        ChannelMessage t;
        t <- mod_3630.get(0);
        mod_3628.put(0, t);
    endrule
    rule rule_4702;
        ChannelMessage t;
        t <- mod_3641.get(0);
        mod_3640.put(1, t);
    endrule
    rule rule_4703;
        ChannelMessage t;
        t <- mod_3626.get(0);
        mod_3626.put(1, t);
    endrule
    rule rule_4704;
        ChannelMessage t;
        t <- mod_3636.get(0);
        mod_3637.put(0, t);
    endrule
    rule rule_4705;
        ChannelMessage t;
        t <- mod_3622.get(0);
        mod_3623.put(0, t);
    endrule
    rule rule_4706;
        ChannelMessage t;
        t <- mod_3648.get(0);
        mod_3648.put(1, t);
    endrule
    rule rule_4707;
        ChannelMessage t;
        t <- mod_3612.get(1);
        mod_3613.put(0, t);
    endrule
    rule rule_4708;
        ChannelMessage t;
        t <- mod_3614.get(1);
        mod_3615.put(0, t);
    endrule
    rule rule_4709;
        ChannelMessage t;
        t <- mod_3612.get(0);
        mod_3648.put(0, t);
    endrule
    rule rule_4710;
        ChannelMessage t;
        t <- mod_3628.get(1);
        mod_3621.put(1, t);
    endrule
    rule rule_4711;
        ChannelMessage t;
        t <- mod_3610.get(0);
        mod_3611.put(0, t);
    endrule
    rule rule_4712;
        ChannelMessage t;
        t <- mod_3611.get(0);
        mod_3612.put(0, t);
    endrule
    rule rule_4713;
        ChannelMessage t;
        t <- mod_3642.get(1);
        mod_3617.put(1, t);
    endrule
    rule rule_4714;
        ChannelMessage t;
        t <- mod_3615.get(0);
        mod_3640.put(0, t);
    endrule
    rule rule_4715;
        ChannelMessage t;
        t <- mod_3627.get(0);
        mod_3627.put(1, t);
    endrule
    rule rule_4716;
        ChannelMessage t;
        t <- mod_3636.get(1);
        mod_3635.put(1, t);
    endrule
    rule rule_4717;
        ChannelMessage t;
        t <- mod_3623.get(0);
        mod_3627.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3609.put(0, t);
        end
        if (i == 1) begin
            mod_3625.put(0, t);
        end
        if (i == 2) begin
            mod_3631.put(0, t);
        end
        if (i == 3) begin
            mod_3639.put(0, t);
        end
        if (i == 4) begin
            mod_3645.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_3613.get(0);
        end
        if (i == 1) begin
            t <- mod_3613.get(1);
        end
        if (i == 0) begin
            t <- mod_3613.get(2);
        end
        if (i == 2) begin
            t <- mod_3625.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6123 (Operation_IFC);
    Operation_IFC mod_3650_inner <- mkReshape(2, 64);
    Operation_IFC mod_3650 <- mkDebugOperation(mod_3650_inner, "mod_3650");
    Operation_IFC mod_3651_inner <- mkFlatten(1);
    Operation_IFC mod_3651 <- mkDebugOperation(mod_3651_inner, "mod_3651");
    Operation_IFC mod_3652_inner <- mkFlatten(2);
    Operation_IFC mod_3652 <- mkDebugOperation(mod_3652_inner, "mod_3652");
    Operation_IFC mod_3653_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3653 <- mkDebugOperation(mod_3653_inner, "mod_3653");
    Broadcast_IFC#(4) mod_3654_inner <- mkBroadcast(4);
    Operation_IFC mod_3654 <- mkDebugOperation(mod_3654_inner.op, "mod_3654");
    PMU_IFC mod_3655_bufferize <- mkPMU(2);
    Operation_IFC mod_3655_inner = mod_3655_bufferize.operation;
    Operation_IFC mod_3655 <- mkDebugOperation(mod_3655_inner, "mod_3655");
    Broadcast_IFC#(2) mod_3656_inner <- mkBroadcast(2);
    Operation_IFC mod_3656 <- mkDebugOperation(mod_3656_inner.op, "mod_3656");
    PMU_IFC mod_3657_bufferize <- mkPMU(1);
    Operation_IFC mod_3657_inner = mod_3657_bufferize.operation;
    Operation_IFC mod_3657 <- mkDebugOperation(mod_3657_inner, "mod_3657");
    Operation_IFC mod_3658_inner <- mkBinaryMap(1067, matmul_t_tile);
    Operation_IFC mod_3658 <- mkDebugOperation(mod_3658_inner, "mod_3658");
    Operation_IFC mod_3659_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3659 <- mkDebugOperation(mod_3659_inner, "mod_3659");
    Operation_IFC mod_3660_inner <- mkBinaryMap(1835, mul_tile);
    Operation_IFC mod_3660 <- mkDebugOperation(mod_3660_inner, "mod_3660");
    PMU_IFC mod_3661_bufferize <- mkPMU(1);
    Operation_IFC mod_3661_inner = mod_3661_bufferize.operation;
    Operation_IFC mod_3661 <- mkDebugOperation(mod_3661_inner, "mod_3661");
    Operation_IFC mod_3662_inner <- mkBinaryMap(2385, matmul_t_tile);
    Operation_IFC mod_3662 <- mkDebugOperation(mod_3662_inner, "mod_3662");
    Operation_IFC mod_3663_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3663 <- mkDebugOperation(mod_3663_inner, "mod_3663");
    Operation_IFC mod_3664_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3664 <- mkDebugOperation(mod_3664_inner, "mod_3664");
    Operation_IFC mod_3665_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3665 <- mkDebugOperation(mod_3665_inner, "mod_3665");
    Operation_IFC mod_3666_inner <- mkBinaryMap(2734, mul_tile);
    Operation_IFC mod_3666 <- mkDebugOperation(mod_3666_inner, "mod_3666");
    PMU_IFC mod_3667_bufferize <- mkPMU(1);
    Operation_IFC mod_3667_inner = mod_3667_bufferize.operation;
    Operation_IFC mod_3667 <- mkDebugOperation(mod_3667_inner, "mod_3667");
    PMU_IFC mod_3668_bufferize <- mkPMU(2);
    Operation_IFC mod_3668_inner = mod_3668_bufferize.operation;
    Operation_IFC mod_3668 <- mkDebugOperation(mod_3668_inner, "mod_3668");
    PMU_IFC mod_3669_bufferize <- mkPMU(2);
    Operation_IFC mod_3669_inner = mod_3669_bufferize.operation;
    Operation_IFC mod_3669 <- mkDebugOperation(mod_3669_inner, "mod_3669");
    Operation_IFC mod_3670_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3670 <- mkDebugOperation(mod_3670_inner, "mod_3670");
    Operation_IFC mod_3671_inner <- mkFlatten(1);
    Operation_IFC mod_3671 <- mkDebugOperation(mod_3671_inner, "mod_3671");
    Operation_IFC mod_3672_inner <- mkFlatten(0);
    Operation_IFC mod_3672 <- mkDebugOperation(mod_3672_inner, "mod_3672");
    Operation_IFC mod_3673_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3673 <- mkDebugOperation(mod_3673_inner, "mod_3673");
    Operation_IFC mod_3674_inner <- mkUnaryMap(1707, silu_tile);
    Operation_IFC mod_3674 <- mkDebugOperation(mod_3674_inner, "mod_3674");
    Operation_IFC mod_3675_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3675 <- mkDebugOperation(mod_3675_inner, "mod_3675");
    Operation_IFC mod_3676_inner <- mkBinaryMap(1579, matmul_t_tile);
    Operation_IFC mod_3676 <- mkDebugOperation(mod_3676_inner, "mod_3676");
    PMU_IFC mod_3677_bufferize <- mkPMU(2);
    Operation_IFC mod_3677_inner = mod_3677_bufferize.operation;
    Operation_IFC mod_3677 <- mkDebugOperation(mod_3677_inner, "mod_3677");
    Operation_IFC mod_3678_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3678 <- mkDebugOperation(mod_3678_inner, "mod_3678");
    Operation_IFC mod_3679_inner <- mkFlatten(1);
    Operation_IFC mod_3679 <- mkDebugOperation(mod_3679_inner, "mod_3679");
    Operation_IFC mod_3680_inner <- mkFlatten(0);
    Operation_IFC mod_3680 <- mkDebugOperation(mod_3680_inner, "mod_3680");
    PMU_IFC mod_3681_bufferize <- mkPMU(1);
    Operation_IFC mod_3681_inner = mod_3681_bufferize.operation;
    Operation_IFC mod_3681 <- mkDebugOperation(mod_3681_inner, "mod_3681");
    Operation_IFC mod_3682_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3682 <- mkDebugOperation(mod_3682_inner, "mod_3682");
    PMU_IFC mod_3683_bufferize <- mkPMU(2);
    Operation_IFC mod_3683_inner = mod_3683_bufferize.operation;
    Operation_IFC mod_3683 <- mkDebugOperation(mod_3683_inner, "mod_3683");
    Operation_IFC mod_3684_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3684 <- mkDebugOperation(mod_3684_inner, "mod_3684");
    Operation_IFC mod_3685_inner <- mkFlatten(1);
    Operation_IFC mod_3685 <- mkDebugOperation(mod_3685_inner, "mod_3685");
    Operation_IFC mod_3686_inner <- mkFlatten(0);
    Operation_IFC mod_3686 <- mkDebugOperation(mod_3686_inner, "mod_3686");
    Operation_IFC mod_3687_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3687 <- mkDebugOperation(mod_3687_inner, "mod_3687");
    Operation_IFC mod_3688_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3688 <- mkDebugOperation(mod_3688_inner, "mod_3688");
    PMU_IFC mod_3689_bufferize <- mkPMU(2);
    Operation_IFC mod_3689_inner = mod_3689_bufferize.operation;
    Operation_IFC mod_3689 <- mkDebugOperation(mod_3689_inner, "mod_3689");
    rule rule_4718;
        ChannelMessage t;
        t <- mod_3681.get(0);
        mod_3682.put(0, t);
    endrule
    rule rule_4719;
        ChannelMessage t;
        t <- mod_3687.get(0);
        mod_3657.put(1, t);
    endrule
    rule rule_4720;
        ChannelMessage t;
        t <- mod_3665.get(0);
        mod_3667.put(0, t);
    endrule
    rule rule_4721;
        ChannelMessage t;
        t <- mod_3664.get(0);
        mod_3668.put(0, t);
    endrule
    rule rule_4722;
        ChannelMessage t;
        t <- mod_3661.get(1);
        mod_3662.put(0, t);
    endrule
    rule rule_4723;
        ChannelMessage t;
        t <- mod_3660.get(0);
        mod_3661.put(0, t);
    endrule
    rule rule_4724;
        ChannelMessage t;
        t <- mod_3689.get(0);
        mod_3689.put(1, t);
    endrule
    rule rule_4725;
        ChannelMessage t;
        t <- mod_3669.get(1);
        mod_3662.put(1, t);
    endrule
    rule rule_4726;
        ChannelMessage t;
        t <- mod_3673.get(0);
        mod_3661.put(1, t);
    endrule
    rule rule_4727;
        ChannelMessage t;
        t <- mod_3670.get(0);
        mod_3669.put(1, t);
    endrule
    rule rule_4728;
        ChannelMessage t;
        t <- mod_3682.get(0);
        mod_3681.put(1, t);
    endrule
    rule rule_4729;
        ChannelMessage t;
        t <- mod_3653.get(0);
        mod_3689.put(0, t);
    endrule
    rule rule_4730;
        ChannelMessage t;
        t <- mod_3651.get(0);
        mod_3652.put(0, t);
    endrule
    rule rule_4731;
        ChannelMessage t;
        t <- mod_3655.get(0);
        mod_3688.put(0, t);
    endrule
    rule rule_4732;
        ChannelMessage t;
        t <- mod_3678.get(0);
        mod_3677.put(1, t);
    endrule
    rule rule_4733;
        ChannelMessage t;
        t <- mod_3661.get(0);
        mod_3673.put(0, t);
    endrule
    rule rule_4734;
        ChannelMessage t;
        t <- mod_3652.get(0);
        mod_3653.put(0, t);
    endrule
    rule rule_4735;
        ChannelMessage t;
        t <- mod_3654.get(3);
        mod_3655.put(0, t);
    endrule
    rule rule_4736;
        ChannelMessage t;
        t <- mod_3668.get(0);
        mod_3668.put(1, t);
    endrule
    rule rule_4737;
        ChannelMessage t;
        t <- mod_3656.get(0);
        mod_3681.put(0, t);
    endrule
    rule rule_4738;
        ChannelMessage t;
        t <- mod_3650.get(0);
        mod_3651.put(0, t);
    endrule
    rule rule_4739;
        ChannelMessage t;
        t <- mod_3659.get(0);
        mod_3660.put(0, t);
    endrule
    rule rule_4740;
        ChannelMessage t;
        t <- mod_3675.get(0);
        mod_3674.put(0, t);
    endrule
    rule rule_4741;
        ChannelMessage t;
        t <- mod_3664.get(1);
        mod_3665.put(0, t);
    endrule
    rule rule_4742;
        ChannelMessage t;
        t <- mod_3677.get(1);
        mod_3676.put(1, t);
    endrule
    rule rule_4743;
        ChannelMessage t;
        t <- mod_3658.get(0);
        mod_3659.put(0, t);
    endrule
    rule rule_4744;
        ChannelMessage t;
        t <- mod_3683.get(1);
        mod_3658.put(1, t);
    endrule
    rule rule_4745;
        ChannelMessage t;
        t <- mod_3667.get(0);
        mod_3667.put(1, t);
    endrule
    rule rule_4746;
        ChannelMessage t;
        t <- mod_3665.get(1);
        mod_3666.put(1, t);
    endrule
    rule rule_4747;
        ChannelMessage t;
        t <- mod_3674.get(0);
        mod_3660.put(1, t);
    endrule
    rule rule_4748;
        ChannelMessage t;
        t <- mod_3667.get(1);
        mod_3665.put(1, t);
    endrule
    rule rule_4749;
        ChannelMessage t;
        t <- mod_3681.get(1);
        mod_3676.put(0, t);
    endrule
    rule rule_4750;
        ChannelMessage t;
        t <- mod_3676.get(0);
        mod_3675.put(0, t);
    endrule
    rule rule_4751;
        ChannelMessage t;
        t <- mod_3677.get(0);
        mod_3678.put(0, t);
    endrule
    rule rule_4752;
        ChannelMessage t;
        t <- mod_3686.get(0);
        mod_3685.put(0, t);
    endrule
    rule rule_4753;
        ChannelMessage t;
        t <- mod_3657.get(0);
        mod_3687.put(0, t);
    endrule
    rule rule_4754;
        ChannelMessage t;
        t <- mod_3685.get(0);
        mod_3683.put(0, t);
    endrule
    rule rule_4755;
        ChannelMessage t;
        t <- mod_3655.get(1);
        mod_3656.put(0, t);
    endrule
    rule rule_4756;
        ChannelMessage t;
        t <- mod_3688.get(0);
        mod_3655.put(1, t);
    endrule
    rule rule_4757;
        ChannelMessage t;
        t <- mod_3684.get(0);
        mod_3683.put(1, t);
    endrule
    rule rule_4758;
        ChannelMessage t;
        t <- mod_3656.get(1);
        mod_3657.put(0, t);
    endrule
    rule rule_4759;
        ChannelMessage t;
        t <- mod_3668.get(1);
        mod_3664.put(1, t);
    endrule
    rule rule_4760;
        ChannelMessage t;
        t <- mod_3683.get(0);
        mod_3684.put(0, t);
    endrule
    rule rule_4761;
        ChannelMessage t;
        t <- mod_3680.get(0);
        mod_3679.put(0, t);
    endrule
    rule rule_4762;
        ChannelMessage t;
        t <- mod_3657.get(1);
        mod_3658.put(0, t);
    endrule
    rule rule_4763;
        ChannelMessage t;
        t <- mod_3662.get(0);
        mod_3663.put(0, t);
    endrule
    rule rule_4764;
        ChannelMessage t;
        t <- mod_3689.get(1);
        mod_3653.put(1, t);
    endrule
    rule rule_4765;
        ChannelMessage t;
        t <- mod_3672.get(0);
        mod_3671.put(0, t);
    endrule
    rule rule_4766;
        ChannelMessage t;
        t <- mod_3653.get(1);
        mod_3654.put(0, t);
    endrule
    rule rule_4767;
        ChannelMessage t;
        t <- mod_3663.get(0);
        mod_3664.put(0, t);
    endrule
    rule rule_4768;
        ChannelMessage t;
        t <- mod_3679.get(0);
        mod_3677.put(0, t);
    endrule
    rule rule_4769;
        ChannelMessage t;
        t <- mod_3671.get(0);
        mod_3669.put(0, t);
    endrule
    rule rule_4770;
        ChannelMessage t;
        t <- mod_3669.get(0);
        mod_3670.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3650.put(0, t);
        end
        if (i == 1) begin
            mod_3666.put(0, t);
        end
        if (i == 2) begin
            mod_3672.put(0, t);
        end
        if (i == 3) begin
            mod_3680.put(0, t);
        end
        if (i == 4) begin
            mod_3686.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_3654.get(0);
        end
        if (i == 2) begin
            t <- mod_3654.get(1);
        end
        if (i == 0) begin
            t <- mod_3654.get(2);
        end
        if (i == 3) begin
            t <- mod_3666.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6124 (Operation_IFC);
    Operation_IFC mod_3691_inner <- mkReshape(2, 64);
    Operation_IFC mod_3691 <- mkDebugOperation(mod_3691_inner, "mod_3691");
    Operation_IFC mod_3692_inner <- mkFlatten(1);
    Operation_IFC mod_3692 <- mkDebugOperation(mod_3692_inner, "mod_3692");
    Operation_IFC mod_3693_inner <- mkFlatten(2);
    Operation_IFC mod_3693 <- mkDebugOperation(mod_3693_inner, "mod_3693");
    Operation_IFC mod_3694_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3694 <- mkDebugOperation(mod_3694_inner, "mod_3694");
    Broadcast_IFC#(4) mod_3695_inner <- mkBroadcast(4);
    Operation_IFC mod_3695 <- mkDebugOperation(mod_3695_inner.op, "mod_3695");
    PMU_IFC mod_3696_bufferize <- mkPMU(2);
    Operation_IFC mod_3696_inner = mod_3696_bufferize.operation;
    Operation_IFC mod_3696 <- mkDebugOperation(mod_3696_inner, "mod_3696");
    Broadcast_IFC#(2) mod_3697_inner <- mkBroadcast(2);
    Operation_IFC mod_3697 <- mkDebugOperation(mod_3697_inner.op, "mod_3697");
    PMU_IFC mod_3698_bufferize <- mkPMU(1);
    Operation_IFC mod_3698_inner = mod_3698_bufferize.operation;
    Operation_IFC mod_3698 <- mkDebugOperation(mod_3698_inner, "mod_3698");
    Operation_IFC mod_3699_inner <- mkBinaryMap(1066, matmul_t_tile);
    Operation_IFC mod_3699 <- mkDebugOperation(mod_3699_inner, "mod_3699");
    Operation_IFC mod_3700_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3700 <- mkDebugOperation(mod_3700_inner, "mod_3700");
    Operation_IFC mod_3701_inner <- mkBinaryMap(1834, mul_tile);
    Operation_IFC mod_3701 <- mkDebugOperation(mod_3701_inner, "mod_3701");
    PMU_IFC mod_3702_bufferize <- mkPMU(1);
    Operation_IFC mod_3702_inner = mod_3702_bufferize.operation;
    Operation_IFC mod_3702 <- mkDebugOperation(mod_3702_inner, "mod_3702");
    Operation_IFC mod_3703_inner <- mkBinaryMap(2383, matmul_t_tile);
    Operation_IFC mod_3703 <- mkDebugOperation(mod_3703_inner, "mod_3703");
    Operation_IFC mod_3704_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3704 <- mkDebugOperation(mod_3704_inner, "mod_3704");
    Operation_IFC mod_3705_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3705 <- mkDebugOperation(mod_3705_inner, "mod_3705");
    Operation_IFC mod_3706_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3706 <- mkDebugOperation(mod_3706_inner, "mod_3706");
    Operation_IFC mod_3707_inner <- mkBinaryMap(2733, mul_tile);
    Operation_IFC mod_3707 <- mkDebugOperation(mod_3707_inner, "mod_3707");
    PMU_IFC mod_3708_bufferize <- mkPMU(1);
    Operation_IFC mod_3708_inner = mod_3708_bufferize.operation;
    Operation_IFC mod_3708 <- mkDebugOperation(mod_3708_inner, "mod_3708");
    PMU_IFC mod_3709_bufferize <- mkPMU(2);
    Operation_IFC mod_3709_inner = mod_3709_bufferize.operation;
    Operation_IFC mod_3709 <- mkDebugOperation(mod_3709_inner, "mod_3709");
    PMU_IFC mod_3710_bufferize <- mkPMU(2);
    Operation_IFC mod_3710_inner = mod_3710_bufferize.operation;
    Operation_IFC mod_3710 <- mkDebugOperation(mod_3710_inner, "mod_3710");
    Operation_IFC mod_3711_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3711 <- mkDebugOperation(mod_3711_inner, "mod_3711");
    Operation_IFC mod_3712_inner <- mkFlatten(1);
    Operation_IFC mod_3712 <- mkDebugOperation(mod_3712_inner, "mod_3712");
    Operation_IFC mod_3713_inner <- mkFlatten(0);
    Operation_IFC mod_3713 <- mkDebugOperation(mod_3713_inner, "mod_3713");
    Operation_IFC mod_3714_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3714 <- mkDebugOperation(mod_3714_inner, "mod_3714");
    Operation_IFC mod_3715_inner <- mkUnaryMap(1706, silu_tile);
    Operation_IFC mod_3715 <- mkDebugOperation(mod_3715_inner, "mod_3715");
    Operation_IFC mod_3716_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3716 <- mkDebugOperation(mod_3716_inner, "mod_3716");
    Operation_IFC mod_3717_inner <- mkBinaryMap(1578, matmul_t_tile);
    Operation_IFC mod_3717 <- mkDebugOperation(mod_3717_inner, "mod_3717");
    PMU_IFC mod_3718_bufferize <- mkPMU(2);
    Operation_IFC mod_3718_inner = mod_3718_bufferize.operation;
    Operation_IFC mod_3718 <- mkDebugOperation(mod_3718_inner, "mod_3718");
    Operation_IFC mod_3719_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3719 <- mkDebugOperation(mod_3719_inner, "mod_3719");
    Operation_IFC mod_3720_inner <- mkFlatten(1);
    Operation_IFC mod_3720 <- mkDebugOperation(mod_3720_inner, "mod_3720");
    Operation_IFC mod_3721_inner <- mkFlatten(0);
    Operation_IFC mod_3721 <- mkDebugOperation(mod_3721_inner, "mod_3721");
    PMU_IFC mod_3722_bufferize <- mkPMU(1);
    Operation_IFC mod_3722_inner = mod_3722_bufferize.operation;
    Operation_IFC mod_3722 <- mkDebugOperation(mod_3722_inner, "mod_3722");
    Operation_IFC mod_3723_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3723 <- mkDebugOperation(mod_3723_inner, "mod_3723");
    PMU_IFC mod_3724_bufferize <- mkPMU(2);
    Operation_IFC mod_3724_inner = mod_3724_bufferize.operation;
    Operation_IFC mod_3724 <- mkDebugOperation(mod_3724_inner, "mod_3724");
    Operation_IFC mod_3725_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3725 <- mkDebugOperation(mod_3725_inner, "mod_3725");
    Operation_IFC mod_3726_inner <- mkFlatten(1);
    Operation_IFC mod_3726 <- mkDebugOperation(mod_3726_inner, "mod_3726");
    Operation_IFC mod_3727_inner <- mkFlatten(0);
    Operation_IFC mod_3727 <- mkDebugOperation(mod_3727_inner, "mod_3727");
    Operation_IFC mod_3728_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3728 <- mkDebugOperation(mod_3728_inner, "mod_3728");
    Operation_IFC mod_3729_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3729 <- mkDebugOperation(mod_3729_inner, "mod_3729");
    PMU_IFC mod_3730_bufferize <- mkPMU(2);
    Operation_IFC mod_3730_inner = mod_3730_bufferize.operation;
    Operation_IFC mod_3730 <- mkDebugOperation(mod_3730_inner, "mod_3730");
    rule rule_4771;
        ChannelMessage t;
        t <- mod_3699.get(0);
        mod_3700.put(0, t);
    endrule
    rule rule_4772;
        ChannelMessage t;
        t <- mod_3712.get(0);
        mod_3710.put(0, t);
    endrule
    rule rule_4773;
        ChannelMessage t;
        t <- mod_3717.get(0);
        mod_3716.put(0, t);
    endrule
    rule rule_4774;
        ChannelMessage t;
        t <- mod_3710.get(0);
        mod_3711.put(0, t);
    endrule
    rule rule_4775;
        ChannelMessage t;
        t <- mod_3692.get(0);
        mod_3693.put(0, t);
    endrule
    rule rule_4776;
        ChannelMessage t;
        t <- mod_3724.get(1);
        mod_3699.put(1, t);
    endrule
    rule rule_4777;
        ChannelMessage t;
        t <- mod_3697.get(1);
        mod_3698.put(0, t);
    endrule
    rule rule_4778;
        ChannelMessage t;
        t <- mod_3695.get(3);
        mod_3696.put(0, t);
    endrule
    rule rule_4779;
        ChannelMessage t;
        t <- mod_3703.get(0);
        mod_3704.put(0, t);
    endrule
    rule rule_4780;
        ChannelMessage t;
        t <- mod_3727.get(0);
        mod_3726.put(0, t);
    endrule
    rule rule_4781;
        ChannelMessage t;
        t <- mod_3706.get(1);
        mod_3707.put(1, t);
    endrule
    rule rule_4782;
        ChannelMessage t;
        t <- mod_3720.get(0);
        mod_3718.put(0, t);
    endrule
    rule rule_4783;
        ChannelMessage t;
        t <- mod_3693.get(0);
        mod_3694.put(0, t);
    endrule
    rule rule_4784;
        ChannelMessage t;
        t <- mod_3730.get(0);
        mod_3730.put(1, t);
    endrule
    rule rule_4785;
        ChannelMessage t;
        t <- mod_3696.get(0);
        mod_3729.put(0, t);
    endrule
    rule rule_4786;
        ChannelMessage t;
        t <- mod_3702.get(1);
        mod_3703.put(0, t);
    endrule
    rule rule_4787;
        ChannelMessage t;
        t <- mod_3723.get(0);
        mod_3722.put(1, t);
    endrule
    rule rule_4788;
        ChannelMessage t;
        t <- mod_3696.get(1);
        mod_3697.put(0, t);
    endrule
    rule rule_4789;
        ChannelMessage t;
        t <- mod_3729.get(0);
        mod_3696.put(1, t);
    endrule
    rule rule_4790;
        ChannelMessage t;
        t <- mod_3704.get(0);
        mod_3705.put(0, t);
    endrule
    rule rule_4791;
        ChannelMessage t;
        t <- mod_3719.get(0);
        mod_3718.put(1, t);
    endrule
    rule rule_4792;
        ChannelMessage t;
        t <- mod_3708.get(1);
        mod_3706.put(1, t);
    endrule
    rule rule_4793;
        ChannelMessage t;
        t <- mod_3691.get(0);
        mod_3692.put(0, t);
    endrule
    rule rule_4794;
        ChannelMessage t;
        t <- mod_3711.get(0);
        mod_3710.put(1, t);
    endrule
    rule rule_4795;
        ChannelMessage t;
        t <- mod_3715.get(0);
        mod_3701.put(1, t);
    endrule
    rule rule_4796;
        ChannelMessage t;
        t <- mod_3700.get(0);
        mod_3701.put(0, t);
    endrule
    rule rule_4797;
        ChannelMessage t;
        t <- mod_3728.get(0);
        mod_3698.put(1, t);
    endrule
    rule rule_4798;
        ChannelMessage t;
        t <- mod_3730.get(1);
        mod_3694.put(1, t);
    endrule
    rule rule_4799;
        ChannelMessage t;
        t <- mod_3706.get(0);
        mod_3708.put(0, t);
    endrule
    rule rule_4800;
        ChannelMessage t;
        t <- mod_3714.get(0);
        mod_3702.put(1, t);
    endrule
    rule rule_4801;
        ChannelMessage t;
        t <- mod_3697.get(0);
        mod_3722.put(0, t);
    endrule
    rule rule_4802;
        ChannelMessage t;
        t <- mod_3716.get(0);
        mod_3715.put(0, t);
    endrule
    rule rule_4803;
        ChannelMessage t;
        t <- mod_3698.get(0);
        mod_3728.put(0, t);
    endrule
    rule rule_4804;
        ChannelMessage t;
        t <- mod_3698.get(1);
        mod_3699.put(0, t);
    endrule
    rule rule_4805;
        ChannelMessage t;
        t <- mod_3694.get(0);
        mod_3730.put(0, t);
    endrule
    rule rule_4806;
        ChannelMessage t;
        t <- mod_3702.get(0);
        mod_3714.put(0, t);
    endrule
    rule rule_4807;
        ChannelMessage t;
        t <- mod_3709.get(0);
        mod_3709.put(1, t);
    endrule
    rule rule_4808;
        ChannelMessage t;
        t <- mod_3721.get(0);
        mod_3720.put(0, t);
    endrule
    rule rule_4809;
        ChannelMessage t;
        t <- mod_3726.get(0);
        mod_3724.put(0, t);
    endrule
    rule rule_4810;
        ChannelMessage t;
        t <- mod_3722.get(0);
        mod_3723.put(0, t);
    endrule
    rule rule_4811;
        ChannelMessage t;
        t <- mod_3701.get(0);
        mod_3702.put(0, t);
    endrule
    rule rule_4812;
        ChannelMessage t;
        t <- mod_3708.get(0);
        mod_3708.put(1, t);
    endrule
    rule rule_4813;
        ChannelMessage t;
        t <- mod_3718.get(1);
        mod_3717.put(1, t);
    endrule
    rule rule_4814;
        ChannelMessage t;
        t <- mod_3713.get(0);
        mod_3712.put(0, t);
    endrule
    rule rule_4815;
        ChannelMessage t;
        t <- mod_3718.get(0);
        mod_3719.put(0, t);
    endrule
    rule rule_4816;
        ChannelMessage t;
        t <- mod_3710.get(1);
        mod_3703.put(1, t);
    endrule
    rule rule_4817;
        ChannelMessage t;
        t <- mod_3725.get(0);
        mod_3724.put(1, t);
    endrule
    rule rule_4818;
        ChannelMessage t;
        t <- mod_3694.get(1);
        mod_3695.put(0, t);
    endrule
    rule rule_4819;
        ChannelMessage t;
        t <- mod_3705.get(1);
        mod_3706.put(0, t);
    endrule
    rule rule_4820;
        ChannelMessage t;
        t <- mod_3705.get(0);
        mod_3709.put(0, t);
    endrule
    rule rule_4821;
        ChannelMessage t;
        t <- mod_3722.get(1);
        mod_3717.put(0, t);
    endrule
    rule rule_4822;
        ChannelMessage t;
        t <- mod_3724.get(0);
        mod_3725.put(0, t);
    endrule
    rule rule_4823;
        ChannelMessage t;
        t <- mod_3709.get(1);
        mod_3705.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3691.put(0, t);
        end
        if (i == 1) begin
            mod_3707.put(0, t);
        end
        if (i == 2) begin
            mod_3713.put(0, t);
        end
        if (i == 3) begin
            mod_3721.put(0, t);
        end
        if (i == 4) begin
            mod_3727.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 2) begin
            t <- mod_3695.get(0);
        end
        if (i == 3) begin
            t <- mod_3695.get(1);
        end
        if (i == 1) begin
            t <- mod_3695.get(2);
        end
        if (i == 0) begin
            t <- mod_3707.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6125 (Operation_IFC);
    Operation_IFC mod_3732_inner <- mkReshape(2, 64);
    Operation_IFC mod_3732 <- mkDebugOperation(mod_3732_inner, "mod_3732");
    Operation_IFC mod_3733_inner <- mkFlatten(1);
    Operation_IFC mod_3733 <- mkDebugOperation(mod_3733_inner, "mod_3733");
    Operation_IFC mod_3734_inner <- mkFlatten(2);
    Operation_IFC mod_3734 <- mkDebugOperation(mod_3734_inner, "mod_3734");
    Operation_IFC mod_3735_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3735 <- mkDebugOperation(mod_3735_inner, "mod_3735");
    Broadcast_IFC#(4) mod_3736_inner <- mkBroadcast(4);
    Operation_IFC mod_3736 <- mkDebugOperation(mod_3736_inner.op, "mod_3736");
    PMU_IFC mod_3737_bufferize <- mkPMU(2);
    Operation_IFC mod_3737_inner = mod_3737_bufferize.operation;
    Operation_IFC mod_3737 <- mkDebugOperation(mod_3737_inner, "mod_3737");
    Broadcast_IFC#(2) mod_3738_inner <- mkBroadcast(2);
    Operation_IFC mod_3738 <- mkDebugOperation(mod_3738_inner.op, "mod_3738");
    PMU_IFC mod_3739_bufferize <- mkPMU(1);
    Operation_IFC mod_3739_inner = mod_3739_bufferize.operation;
    Operation_IFC mod_3739 <- mkDebugOperation(mod_3739_inner, "mod_3739");
    Operation_IFC mod_3740_inner <- mkBinaryMap(1065, matmul_t_tile);
    Operation_IFC mod_3740 <- mkDebugOperation(mod_3740_inner, "mod_3740");
    Operation_IFC mod_3741_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3741 <- mkDebugOperation(mod_3741_inner, "mod_3741");
    Operation_IFC mod_3742_inner <- mkBinaryMap(1833, mul_tile);
    Operation_IFC mod_3742 <- mkDebugOperation(mod_3742_inner, "mod_3742");
    PMU_IFC mod_3743_bufferize <- mkPMU(1);
    Operation_IFC mod_3743_inner = mod_3743_bufferize.operation;
    Operation_IFC mod_3743 <- mkDebugOperation(mod_3743_inner, "mod_3743");
    Operation_IFC mod_3744_inner <- mkBinaryMap(2381, matmul_t_tile);
    Operation_IFC mod_3744 <- mkDebugOperation(mod_3744_inner, "mod_3744");
    Operation_IFC mod_3745_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3745 <- mkDebugOperation(mod_3745_inner, "mod_3745");
    Operation_IFC mod_3746_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3746 <- mkDebugOperation(mod_3746_inner, "mod_3746");
    Operation_IFC mod_3747_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3747 <- mkDebugOperation(mod_3747_inner, "mod_3747");
    Operation_IFC mod_3748_inner <- mkBinaryMap(2732, mul_tile);
    Operation_IFC mod_3748 <- mkDebugOperation(mod_3748_inner, "mod_3748");
    PMU_IFC mod_3749_bufferize <- mkPMU(1);
    Operation_IFC mod_3749_inner = mod_3749_bufferize.operation;
    Operation_IFC mod_3749 <- mkDebugOperation(mod_3749_inner, "mod_3749");
    PMU_IFC mod_3750_bufferize <- mkPMU(2);
    Operation_IFC mod_3750_inner = mod_3750_bufferize.operation;
    Operation_IFC mod_3750 <- mkDebugOperation(mod_3750_inner, "mod_3750");
    PMU_IFC mod_3751_bufferize <- mkPMU(2);
    Operation_IFC mod_3751_inner = mod_3751_bufferize.operation;
    Operation_IFC mod_3751 <- mkDebugOperation(mod_3751_inner, "mod_3751");
    Operation_IFC mod_3752_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3752 <- mkDebugOperation(mod_3752_inner, "mod_3752");
    Operation_IFC mod_3753_inner <- mkFlatten(1);
    Operation_IFC mod_3753 <- mkDebugOperation(mod_3753_inner, "mod_3753");
    Operation_IFC mod_3754_inner <- mkFlatten(0);
    Operation_IFC mod_3754 <- mkDebugOperation(mod_3754_inner, "mod_3754");
    Operation_IFC mod_3755_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3755 <- mkDebugOperation(mod_3755_inner, "mod_3755");
    Operation_IFC mod_3756_inner <- mkUnaryMap(1705, silu_tile);
    Operation_IFC mod_3756 <- mkDebugOperation(mod_3756_inner, "mod_3756");
    Operation_IFC mod_3757_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3757 <- mkDebugOperation(mod_3757_inner, "mod_3757");
    Operation_IFC mod_3758_inner <- mkBinaryMap(1577, matmul_t_tile);
    Operation_IFC mod_3758 <- mkDebugOperation(mod_3758_inner, "mod_3758");
    PMU_IFC mod_3759_bufferize <- mkPMU(2);
    Operation_IFC mod_3759_inner = mod_3759_bufferize.operation;
    Operation_IFC mod_3759 <- mkDebugOperation(mod_3759_inner, "mod_3759");
    Operation_IFC mod_3760_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3760 <- mkDebugOperation(mod_3760_inner, "mod_3760");
    Operation_IFC mod_3761_inner <- mkFlatten(1);
    Operation_IFC mod_3761 <- mkDebugOperation(mod_3761_inner, "mod_3761");
    Operation_IFC mod_3762_inner <- mkFlatten(0);
    Operation_IFC mod_3762 <- mkDebugOperation(mod_3762_inner, "mod_3762");
    PMU_IFC mod_3763_bufferize <- mkPMU(1);
    Operation_IFC mod_3763_inner = mod_3763_bufferize.operation;
    Operation_IFC mod_3763 <- mkDebugOperation(mod_3763_inner, "mod_3763");
    Operation_IFC mod_3764_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3764 <- mkDebugOperation(mod_3764_inner, "mod_3764");
    PMU_IFC mod_3765_bufferize <- mkPMU(2);
    Operation_IFC mod_3765_inner = mod_3765_bufferize.operation;
    Operation_IFC mod_3765 <- mkDebugOperation(mod_3765_inner, "mod_3765");
    Operation_IFC mod_3766_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3766 <- mkDebugOperation(mod_3766_inner, "mod_3766");
    Operation_IFC mod_3767_inner <- mkFlatten(1);
    Operation_IFC mod_3767 <- mkDebugOperation(mod_3767_inner, "mod_3767");
    Operation_IFC mod_3768_inner <- mkFlatten(0);
    Operation_IFC mod_3768 <- mkDebugOperation(mod_3768_inner, "mod_3768");
    Operation_IFC mod_3769_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3769 <- mkDebugOperation(mod_3769_inner, "mod_3769");
    Operation_IFC mod_3770_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3770 <- mkDebugOperation(mod_3770_inner, "mod_3770");
    PMU_IFC mod_3771_bufferize <- mkPMU(2);
    Operation_IFC mod_3771_inner = mod_3771_bufferize.operation;
    Operation_IFC mod_3771 <- mkDebugOperation(mod_3771_inner, "mod_3771");
    rule rule_4824;
        ChannelMessage t;
        t <- mod_3765.get(0);
        mod_3766.put(0, t);
    endrule
    rule rule_4825;
        ChannelMessage t;
        t <- mod_3737.get(1);
        mod_3738.put(0, t);
    endrule
    rule rule_4826;
        ChannelMessage t;
        t <- mod_3734.get(0);
        mod_3735.put(0, t);
    endrule
    rule rule_4827;
        ChannelMessage t;
        t <- mod_3764.get(0);
        mod_3763.put(1, t);
    endrule
    rule rule_4828;
        ChannelMessage t;
        t <- mod_3747.get(1);
        mod_3748.put(1, t);
    endrule
    rule rule_4829;
        ChannelMessage t;
        t <- mod_3766.get(0);
        mod_3765.put(1, t);
    endrule
    rule rule_4830;
        ChannelMessage t;
        t <- mod_3771.get(1);
        mod_3735.put(1, t);
    endrule
    rule rule_4831;
        ChannelMessage t;
        t <- mod_3743.get(1);
        mod_3744.put(0, t);
    endrule
    rule rule_4832;
        ChannelMessage t;
        t <- mod_3751.get(1);
        mod_3744.put(1, t);
    endrule
    rule rule_4833;
        ChannelMessage t;
        t <- mod_3749.get(0);
        mod_3749.put(1, t);
    endrule
    rule rule_4834;
        ChannelMessage t;
        t <- mod_3746.get(0);
        mod_3750.put(0, t);
    endrule
    rule rule_4835;
        ChannelMessage t;
        t <- mod_3758.get(0);
        mod_3757.put(0, t);
    endrule
    rule rule_4836;
        ChannelMessage t;
        t <- mod_3750.get(1);
        mod_3746.put(1, t);
    endrule
    rule rule_4837;
        ChannelMessage t;
        t <- mod_3737.get(0);
        mod_3770.put(0, t);
    endrule
    rule rule_4838;
        ChannelMessage t;
        t <- mod_3740.get(0);
        mod_3741.put(0, t);
    endrule
    rule rule_4839;
        ChannelMessage t;
        t <- mod_3732.get(0);
        mod_3733.put(0, t);
    endrule
    rule rule_4840;
        ChannelMessage t;
        t <- mod_3754.get(0);
        mod_3753.put(0, t);
    endrule
    rule rule_4841;
        ChannelMessage t;
        t <- mod_3759.get(0);
        mod_3760.put(0, t);
    endrule
    rule rule_4842;
        ChannelMessage t;
        t <- mod_3743.get(0);
        mod_3755.put(0, t);
    endrule
    rule rule_4843;
        ChannelMessage t;
        t <- mod_3744.get(0);
        mod_3745.put(0, t);
    endrule
    rule rule_4844;
        ChannelMessage t;
        t <- mod_3739.get(1);
        mod_3740.put(0, t);
    endrule
    rule rule_4845;
        ChannelMessage t;
        t <- mod_3763.get(1);
        mod_3758.put(0, t);
    endrule
    rule rule_4846;
        ChannelMessage t;
        t <- mod_3738.get(0);
        mod_3763.put(0, t);
    endrule
    rule rule_4847;
        ChannelMessage t;
        t <- mod_3767.get(0);
        mod_3765.put(0, t);
    endrule
    rule rule_4848;
        ChannelMessage t;
        t <- mod_3761.get(0);
        mod_3759.put(0, t);
    endrule
    rule rule_4849;
        ChannelMessage t;
        t <- mod_3768.get(0);
        mod_3767.put(0, t);
    endrule
    rule rule_4850;
        ChannelMessage t;
        t <- mod_3769.get(0);
        mod_3739.put(1, t);
    endrule
    rule rule_4851;
        ChannelMessage t;
        t <- mod_3735.get(0);
        mod_3771.put(0, t);
    endrule
    rule rule_4852;
        ChannelMessage t;
        t <- mod_3750.get(0);
        mod_3750.put(1, t);
    endrule
    rule rule_4853;
        ChannelMessage t;
        t <- mod_3771.get(0);
        mod_3771.put(1, t);
    endrule
    rule rule_4854;
        ChannelMessage t;
        t <- mod_3757.get(0);
        mod_3756.put(0, t);
    endrule
    rule rule_4855;
        ChannelMessage t;
        t <- mod_3733.get(0);
        mod_3734.put(0, t);
    endrule
    rule rule_4856;
        ChannelMessage t;
        t <- mod_3763.get(0);
        mod_3764.put(0, t);
    endrule
    rule rule_4857;
        ChannelMessage t;
        t <- mod_3751.get(0);
        mod_3752.put(0, t);
    endrule
    rule rule_4858;
        ChannelMessage t;
        t <- mod_3749.get(1);
        mod_3747.put(1, t);
    endrule
    rule rule_4859;
        ChannelMessage t;
        t <- mod_3755.get(0);
        mod_3743.put(1, t);
    endrule
    rule rule_4860;
        ChannelMessage t;
        t <- mod_3741.get(0);
        mod_3742.put(0, t);
    endrule
    rule rule_4861;
        ChannelMessage t;
        t <- mod_3747.get(0);
        mod_3749.put(0, t);
    endrule
    rule rule_4862;
        ChannelMessage t;
        t <- mod_3735.get(1);
        mod_3736.put(0, t);
    endrule
    rule rule_4863;
        ChannelMessage t;
        t <- mod_3759.get(1);
        mod_3758.put(1, t);
    endrule
    rule rule_4864;
        ChannelMessage t;
        t <- mod_3765.get(1);
        mod_3740.put(1, t);
    endrule
    rule rule_4865;
        ChannelMessage t;
        t <- mod_3738.get(1);
        mod_3739.put(0, t);
    endrule
    rule rule_4866;
        ChannelMessage t;
        t <- mod_3756.get(0);
        mod_3742.put(1, t);
    endrule
    rule rule_4867;
        ChannelMessage t;
        t <- mod_3745.get(0);
        mod_3746.put(0, t);
    endrule
    rule rule_4868;
        ChannelMessage t;
        t <- mod_3760.get(0);
        mod_3759.put(1, t);
    endrule
    rule rule_4869;
        ChannelMessage t;
        t <- mod_3762.get(0);
        mod_3761.put(0, t);
    endrule
    rule rule_4870;
        ChannelMessage t;
        t <- mod_3770.get(0);
        mod_3737.put(1, t);
    endrule
    rule rule_4871;
        ChannelMessage t;
        t <- mod_3742.get(0);
        mod_3743.put(0, t);
    endrule
    rule rule_4872;
        ChannelMessage t;
        t <- mod_3746.get(1);
        mod_3747.put(0, t);
    endrule
    rule rule_4873;
        ChannelMessage t;
        t <- mod_3736.get(3);
        mod_3737.put(0, t);
    endrule
    rule rule_4874;
        ChannelMessage t;
        t <- mod_3752.get(0);
        mod_3751.put(1, t);
    endrule
    rule rule_4875;
        ChannelMessage t;
        t <- mod_3753.get(0);
        mod_3751.put(0, t);
    endrule
    rule rule_4876;
        ChannelMessage t;
        t <- mod_3739.get(0);
        mod_3769.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3732.put(0, t);
        end
        if (i == 1) begin
            mod_3748.put(0, t);
        end
        if (i == 2) begin
            mod_3754.put(0, t);
        end
        if (i == 3) begin
            mod_3762.put(0, t);
        end
        if (i == 4) begin
            mod_3768.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 2) begin
            t <- mod_3736.get(0);
        end
        if (i == 0) begin
            t <- mod_3736.get(1);
        end
        if (i == 3) begin
            t <- mod_3736.get(2);
        end
        if (i == 1) begin
            t <- mod_3748.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6126 (Operation_IFC);
    Operation_IFC mod_3773_inner <- mkReshape(2, 64);
    Operation_IFC mod_3773 <- mkDebugOperation(mod_3773_inner, "mod_3773");
    Operation_IFC mod_3774_inner <- mkFlatten(1);
    Operation_IFC mod_3774 <- mkDebugOperation(mod_3774_inner, "mod_3774");
    Operation_IFC mod_3775_inner <- mkFlatten(2);
    Operation_IFC mod_3775 <- mkDebugOperation(mod_3775_inner, "mod_3775");
    Operation_IFC mod_3776_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3776 <- mkDebugOperation(mod_3776_inner, "mod_3776");
    Broadcast_IFC#(4) mod_3777_inner <- mkBroadcast(4);
    Operation_IFC mod_3777 <- mkDebugOperation(mod_3777_inner.op, "mod_3777");
    PMU_IFC mod_3778_bufferize <- mkPMU(2);
    Operation_IFC mod_3778_inner = mod_3778_bufferize.operation;
    Operation_IFC mod_3778 <- mkDebugOperation(mod_3778_inner, "mod_3778");
    Broadcast_IFC#(2) mod_3779_inner <- mkBroadcast(2);
    Operation_IFC mod_3779 <- mkDebugOperation(mod_3779_inner.op, "mod_3779");
    PMU_IFC mod_3780_bufferize <- mkPMU(1);
    Operation_IFC mod_3780_inner = mod_3780_bufferize.operation;
    Operation_IFC mod_3780 <- mkDebugOperation(mod_3780_inner, "mod_3780");
    Operation_IFC mod_3781_inner <- mkBinaryMap(1064, matmul_t_tile);
    Operation_IFC mod_3781 <- mkDebugOperation(mod_3781_inner, "mod_3781");
    Operation_IFC mod_3782_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3782 <- mkDebugOperation(mod_3782_inner, "mod_3782");
    Operation_IFC mod_3783_inner <- mkBinaryMap(1832, mul_tile);
    Operation_IFC mod_3783 <- mkDebugOperation(mod_3783_inner, "mod_3783");
    PMU_IFC mod_3784_bufferize <- mkPMU(1);
    Operation_IFC mod_3784_inner = mod_3784_bufferize.operation;
    Operation_IFC mod_3784 <- mkDebugOperation(mod_3784_inner, "mod_3784");
    Operation_IFC mod_3785_inner <- mkBinaryMap(2379, matmul_t_tile);
    Operation_IFC mod_3785 <- mkDebugOperation(mod_3785_inner, "mod_3785");
    Operation_IFC mod_3786_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3786 <- mkDebugOperation(mod_3786_inner, "mod_3786");
    Operation_IFC mod_3787_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3787 <- mkDebugOperation(mod_3787_inner, "mod_3787");
    Operation_IFC mod_3788_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3788 <- mkDebugOperation(mod_3788_inner, "mod_3788");
    Operation_IFC mod_3789_inner <- mkBinaryMap(2731, mul_tile);
    Operation_IFC mod_3789 <- mkDebugOperation(mod_3789_inner, "mod_3789");
    PMU_IFC mod_3790_bufferize <- mkPMU(1);
    Operation_IFC mod_3790_inner = mod_3790_bufferize.operation;
    Operation_IFC mod_3790 <- mkDebugOperation(mod_3790_inner, "mod_3790");
    PMU_IFC mod_3791_bufferize <- mkPMU(2);
    Operation_IFC mod_3791_inner = mod_3791_bufferize.operation;
    Operation_IFC mod_3791 <- mkDebugOperation(mod_3791_inner, "mod_3791");
    PMU_IFC mod_3792_bufferize <- mkPMU(2);
    Operation_IFC mod_3792_inner = mod_3792_bufferize.operation;
    Operation_IFC mod_3792 <- mkDebugOperation(mod_3792_inner, "mod_3792");
    Operation_IFC mod_3793_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3793 <- mkDebugOperation(mod_3793_inner, "mod_3793");
    Operation_IFC mod_3794_inner <- mkFlatten(1);
    Operation_IFC mod_3794 <- mkDebugOperation(mod_3794_inner, "mod_3794");
    Operation_IFC mod_3795_inner <- mkFlatten(0);
    Operation_IFC mod_3795 <- mkDebugOperation(mod_3795_inner, "mod_3795");
    Operation_IFC mod_3796_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3796 <- mkDebugOperation(mod_3796_inner, "mod_3796");
    Operation_IFC mod_3797_inner <- mkUnaryMap(1704, silu_tile);
    Operation_IFC mod_3797 <- mkDebugOperation(mod_3797_inner, "mod_3797");
    Operation_IFC mod_3798_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3798 <- mkDebugOperation(mod_3798_inner, "mod_3798");
    Operation_IFC mod_3799_inner <- mkBinaryMap(1576, matmul_t_tile);
    Operation_IFC mod_3799 <- mkDebugOperation(mod_3799_inner, "mod_3799");
    PMU_IFC mod_3800_bufferize <- mkPMU(2);
    Operation_IFC mod_3800_inner = mod_3800_bufferize.operation;
    Operation_IFC mod_3800 <- mkDebugOperation(mod_3800_inner, "mod_3800");
    Operation_IFC mod_3801_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3801 <- mkDebugOperation(mod_3801_inner, "mod_3801");
    Operation_IFC mod_3802_inner <- mkFlatten(1);
    Operation_IFC mod_3802 <- mkDebugOperation(mod_3802_inner, "mod_3802");
    Operation_IFC mod_3803_inner <- mkFlatten(0);
    Operation_IFC mod_3803 <- mkDebugOperation(mod_3803_inner, "mod_3803");
    PMU_IFC mod_3804_bufferize <- mkPMU(1);
    Operation_IFC mod_3804_inner = mod_3804_bufferize.operation;
    Operation_IFC mod_3804 <- mkDebugOperation(mod_3804_inner, "mod_3804");
    Operation_IFC mod_3805_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3805 <- mkDebugOperation(mod_3805_inner, "mod_3805");
    PMU_IFC mod_3806_bufferize <- mkPMU(2);
    Operation_IFC mod_3806_inner = mod_3806_bufferize.operation;
    Operation_IFC mod_3806 <- mkDebugOperation(mod_3806_inner, "mod_3806");
    Operation_IFC mod_3807_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3807 <- mkDebugOperation(mod_3807_inner, "mod_3807");
    Operation_IFC mod_3808_inner <- mkFlatten(1);
    Operation_IFC mod_3808 <- mkDebugOperation(mod_3808_inner, "mod_3808");
    Operation_IFC mod_3809_inner <- mkFlatten(0);
    Operation_IFC mod_3809 <- mkDebugOperation(mod_3809_inner, "mod_3809");
    Operation_IFC mod_3810_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3810 <- mkDebugOperation(mod_3810_inner, "mod_3810");
    Operation_IFC mod_3811_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3811 <- mkDebugOperation(mod_3811_inner, "mod_3811");
    PMU_IFC mod_3812_bufferize <- mkPMU(2);
    Operation_IFC mod_3812_inner = mod_3812_bufferize.operation;
    Operation_IFC mod_3812 <- mkDebugOperation(mod_3812_inner, "mod_3812");
    rule rule_4877;
        ChannelMessage t;
        t <- mod_3797.get(0);
        mod_3783.put(1, t);
    endrule
    rule rule_4878;
        ChannelMessage t;
        t <- mod_3795.get(0);
        mod_3794.put(0, t);
    endrule
    rule rule_4879;
        ChannelMessage t;
        t <- mod_3775.get(0);
        mod_3776.put(0, t);
    endrule
    rule rule_4880;
        ChannelMessage t;
        t <- mod_3776.get(1);
        mod_3777.put(0, t);
    endrule
    rule rule_4881;
        ChannelMessage t;
        t <- mod_3785.get(0);
        mod_3786.put(0, t);
    endrule
    rule rule_4882;
        ChannelMessage t;
        t <- mod_3804.get(1);
        mod_3799.put(0, t);
    endrule
    rule rule_4883;
        ChannelMessage t;
        t <- mod_3810.get(0);
        mod_3780.put(1, t);
    endrule
    rule rule_4884;
        ChannelMessage t;
        t <- mod_3783.get(0);
        mod_3784.put(0, t);
    endrule
    rule rule_4885;
        ChannelMessage t;
        t <- mod_3807.get(0);
        mod_3806.put(1, t);
    endrule
    rule rule_4886;
        ChannelMessage t;
        t <- mod_3773.get(0);
        mod_3774.put(0, t);
    endrule
    rule rule_4887;
        ChannelMessage t;
        t <- mod_3803.get(0);
        mod_3802.put(0, t);
    endrule
    rule rule_4888;
        ChannelMessage t;
        t <- mod_3806.get(1);
        mod_3781.put(1, t);
    endrule
    rule rule_4889;
        ChannelMessage t;
        t <- mod_3791.get(1);
        mod_3787.put(1, t);
    endrule
    rule rule_4890;
        ChannelMessage t;
        t <- mod_3790.get(0);
        mod_3790.put(1, t);
    endrule
    rule rule_4891;
        ChannelMessage t;
        t <- mod_3805.get(0);
        mod_3804.put(1, t);
    endrule
    rule rule_4892;
        ChannelMessage t;
        t <- mod_3780.get(1);
        mod_3781.put(0, t);
    endrule
    rule rule_4893;
        ChannelMessage t;
        t <- mod_3790.get(1);
        mod_3788.put(1, t);
    endrule
    rule rule_4894;
        ChannelMessage t;
        t <- mod_3801.get(0);
        mod_3800.put(1, t);
    endrule
    rule rule_4895;
        ChannelMessage t;
        t <- mod_3784.get(1);
        mod_3785.put(0, t);
    endrule
    rule rule_4896;
        ChannelMessage t;
        t <- mod_3798.get(0);
        mod_3797.put(0, t);
    endrule
    rule rule_4897;
        ChannelMessage t;
        t <- mod_3778.get(0);
        mod_3811.put(0, t);
    endrule
    rule rule_4898;
        ChannelMessage t;
        t <- mod_3777.get(3);
        mod_3778.put(0, t);
    endrule
    rule rule_4899;
        ChannelMessage t;
        t <- mod_3808.get(0);
        mod_3806.put(0, t);
    endrule
    rule rule_4900;
        ChannelMessage t;
        t <- mod_3774.get(0);
        mod_3775.put(0, t);
    endrule
    rule rule_4901;
        ChannelMessage t;
        t <- mod_3776.get(0);
        mod_3812.put(0, t);
    endrule
    rule rule_4902;
        ChannelMessage t;
        t <- mod_3779.get(0);
        mod_3804.put(0, t);
    endrule
    rule rule_4903;
        ChannelMessage t;
        t <- mod_3782.get(0);
        mod_3783.put(0, t);
    endrule
    rule rule_4904;
        ChannelMessage t;
        t <- mod_3787.get(0);
        mod_3791.put(0, t);
    endrule
    rule rule_4905;
        ChannelMessage t;
        t <- mod_3792.get(1);
        mod_3785.put(1, t);
    endrule
    rule rule_4906;
        ChannelMessage t;
        t <- mod_3800.get(0);
        mod_3801.put(0, t);
    endrule
    rule rule_4907;
        ChannelMessage t;
        t <- mod_3784.get(0);
        mod_3796.put(0, t);
    endrule
    rule rule_4908;
        ChannelMessage t;
        t <- mod_3793.get(0);
        mod_3792.put(1, t);
    endrule
    rule rule_4909;
        ChannelMessage t;
        t <- mod_3812.get(1);
        mod_3776.put(1, t);
    endrule
    rule rule_4910;
        ChannelMessage t;
        t <- mod_3778.get(1);
        mod_3779.put(0, t);
    endrule
    rule rule_4911;
        ChannelMessage t;
        t <- mod_3802.get(0);
        mod_3800.put(0, t);
    endrule
    rule rule_4912;
        ChannelMessage t;
        t <- mod_3781.get(0);
        mod_3782.put(0, t);
    endrule
    rule rule_4913;
        ChannelMessage t;
        t <- mod_3812.get(0);
        mod_3812.put(1, t);
    endrule
    rule rule_4914;
        ChannelMessage t;
        t <- mod_3788.get(0);
        mod_3790.put(0, t);
    endrule
    rule rule_4915;
        ChannelMessage t;
        t <- mod_3788.get(1);
        mod_3789.put(1, t);
    endrule
    rule rule_4916;
        ChannelMessage t;
        t <- mod_3809.get(0);
        mod_3808.put(0, t);
    endrule
    rule rule_4917;
        ChannelMessage t;
        t <- mod_3779.get(1);
        mod_3780.put(0, t);
    endrule
    rule rule_4918;
        ChannelMessage t;
        t <- mod_3780.get(0);
        mod_3810.put(0, t);
    endrule
    rule rule_4919;
        ChannelMessage t;
        t <- mod_3806.get(0);
        mod_3807.put(0, t);
    endrule
    rule rule_4920;
        ChannelMessage t;
        t <- mod_3791.get(0);
        mod_3791.put(1, t);
    endrule
    rule rule_4921;
        ChannelMessage t;
        t <- mod_3792.get(0);
        mod_3793.put(0, t);
    endrule
    rule rule_4922;
        ChannelMessage t;
        t <- mod_3787.get(1);
        mod_3788.put(0, t);
    endrule
    rule rule_4923;
        ChannelMessage t;
        t <- mod_3799.get(0);
        mod_3798.put(0, t);
    endrule
    rule rule_4924;
        ChannelMessage t;
        t <- mod_3786.get(0);
        mod_3787.put(0, t);
    endrule
    rule rule_4925;
        ChannelMessage t;
        t <- mod_3796.get(0);
        mod_3784.put(1, t);
    endrule
    rule rule_4926;
        ChannelMessage t;
        t <- mod_3800.get(1);
        mod_3799.put(1, t);
    endrule
    rule rule_4927;
        ChannelMessage t;
        t <- mod_3811.get(0);
        mod_3778.put(1, t);
    endrule
    rule rule_4928;
        ChannelMessage t;
        t <- mod_3794.get(0);
        mod_3792.put(0, t);
    endrule
    rule rule_4929;
        ChannelMessage t;
        t <- mod_3804.get(0);
        mod_3805.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3773.put(0, t);
        end
        if (i == 1) begin
            mod_3789.put(0, t);
        end
        if (i == 2) begin
            mod_3795.put(0, t);
        end
        if (i == 3) begin
            mod_3803.put(0, t);
        end
        if (i == 4) begin
            mod_3809.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_3777.get(0);
        end
        if (i == 2) begin
            t <- mod_3777.get(1);
        end
        if (i == 3) begin
            t <- mod_3777.get(2);
        end
        if (i == 1) begin
            t <- mod_3789.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6127 (Operation_IFC);
    Operation_IFC mod_3814_inner <- mkReshape(2, 64);
    Operation_IFC mod_3814 <- mkDebugOperation(mod_3814_inner, "mod_3814");
    Operation_IFC mod_3815_inner <- mkFlatten(1);
    Operation_IFC mod_3815 <- mkDebugOperation(mod_3815_inner, "mod_3815");
    Operation_IFC mod_3816_inner <- mkFlatten(2);
    Operation_IFC mod_3816 <- mkDebugOperation(mod_3816_inner, "mod_3816");
    Operation_IFC mod_3817_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3817 <- mkDebugOperation(mod_3817_inner, "mod_3817");
    Broadcast_IFC#(4) mod_3818_inner <- mkBroadcast(4);
    Operation_IFC mod_3818 <- mkDebugOperation(mod_3818_inner.op, "mod_3818");
    PMU_IFC mod_3819_bufferize <- mkPMU(2);
    Operation_IFC mod_3819_inner = mod_3819_bufferize.operation;
    Operation_IFC mod_3819 <- mkDebugOperation(mod_3819_inner, "mod_3819");
    Broadcast_IFC#(2) mod_3820_inner <- mkBroadcast(2);
    Operation_IFC mod_3820 <- mkDebugOperation(mod_3820_inner.op, "mod_3820");
    PMU_IFC mod_3821_bufferize <- mkPMU(1);
    Operation_IFC mod_3821_inner = mod_3821_bufferize.operation;
    Operation_IFC mod_3821 <- mkDebugOperation(mod_3821_inner, "mod_3821");
    Operation_IFC mod_3822_inner <- mkBinaryMap(1063, matmul_t_tile);
    Operation_IFC mod_3822 <- mkDebugOperation(mod_3822_inner, "mod_3822");
    Operation_IFC mod_3823_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3823 <- mkDebugOperation(mod_3823_inner, "mod_3823");
    Operation_IFC mod_3824_inner <- mkBinaryMap(1831, mul_tile);
    Operation_IFC mod_3824 <- mkDebugOperation(mod_3824_inner, "mod_3824");
    PMU_IFC mod_3825_bufferize <- mkPMU(1);
    Operation_IFC mod_3825_inner = mod_3825_bufferize.operation;
    Operation_IFC mod_3825 <- mkDebugOperation(mod_3825_inner, "mod_3825");
    Operation_IFC mod_3826_inner <- mkBinaryMap(2377, matmul_t_tile);
    Operation_IFC mod_3826 <- mkDebugOperation(mod_3826_inner, "mod_3826");
    Operation_IFC mod_3827_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3827 <- mkDebugOperation(mod_3827_inner, "mod_3827");
    Operation_IFC mod_3828_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3828 <- mkDebugOperation(mod_3828_inner, "mod_3828");
    Operation_IFC mod_3829_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3829 <- mkDebugOperation(mod_3829_inner, "mod_3829");
    Operation_IFC mod_3830_inner <- mkBinaryMap(2730, mul_tile);
    Operation_IFC mod_3830 <- mkDebugOperation(mod_3830_inner, "mod_3830");
    PMU_IFC mod_3831_bufferize <- mkPMU(1);
    Operation_IFC mod_3831_inner = mod_3831_bufferize.operation;
    Operation_IFC mod_3831 <- mkDebugOperation(mod_3831_inner, "mod_3831");
    PMU_IFC mod_3832_bufferize <- mkPMU(2);
    Operation_IFC mod_3832_inner = mod_3832_bufferize.operation;
    Operation_IFC mod_3832 <- mkDebugOperation(mod_3832_inner, "mod_3832");
    PMU_IFC mod_3833_bufferize <- mkPMU(2);
    Operation_IFC mod_3833_inner = mod_3833_bufferize.operation;
    Operation_IFC mod_3833 <- mkDebugOperation(mod_3833_inner, "mod_3833");
    Operation_IFC mod_3834_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3834 <- mkDebugOperation(mod_3834_inner, "mod_3834");
    Operation_IFC mod_3835_inner <- mkFlatten(1);
    Operation_IFC mod_3835 <- mkDebugOperation(mod_3835_inner, "mod_3835");
    Operation_IFC mod_3836_inner <- mkFlatten(0);
    Operation_IFC mod_3836 <- mkDebugOperation(mod_3836_inner, "mod_3836");
    Operation_IFC mod_3837_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3837 <- mkDebugOperation(mod_3837_inner, "mod_3837");
    Operation_IFC mod_3838_inner <- mkUnaryMap(1703, silu_tile);
    Operation_IFC mod_3838 <- mkDebugOperation(mod_3838_inner, "mod_3838");
    Operation_IFC mod_3839_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3839 <- mkDebugOperation(mod_3839_inner, "mod_3839");
    Operation_IFC mod_3840_inner <- mkBinaryMap(1575, matmul_t_tile);
    Operation_IFC mod_3840 <- mkDebugOperation(mod_3840_inner, "mod_3840");
    PMU_IFC mod_3841_bufferize <- mkPMU(2);
    Operation_IFC mod_3841_inner = mod_3841_bufferize.operation;
    Operation_IFC mod_3841 <- mkDebugOperation(mod_3841_inner, "mod_3841");
    Operation_IFC mod_3842_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3842 <- mkDebugOperation(mod_3842_inner, "mod_3842");
    Operation_IFC mod_3843_inner <- mkFlatten(1);
    Operation_IFC mod_3843 <- mkDebugOperation(mod_3843_inner, "mod_3843");
    Operation_IFC mod_3844_inner <- mkFlatten(0);
    Operation_IFC mod_3844 <- mkDebugOperation(mod_3844_inner, "mod_3844");
    PMU_IFC mod_3845_bufferize <- mkPMU(1);
    Operation_IFC mod_3845_inner = mod_3845_bufferize.operation;
    Operation_IFC mod_3845 <- mkDebugOperation(mod_3845_inner, "mod_3845");
    Operation_IFC mod_3846_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3846 <- mkDebugOperation(mod_3846_inner, "mod_3846");
    PMU_IFC mod_3847_bufferize <- mkPMU(2);
    Operation_IFC mod_3847_inner = mod_3847_bufferize.operation;
    Operation_IFC mod_3847 <- mkDebugOperation(mod_3847_inner, "mod_3847");
    Operation_IFC mod_3848_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3848 <- mkDebugOperation(mod_3848_inner, "mod_3848");
    Operation_IFC mod_3849_inner <- mkFlatten(1);
    Operation_IFC mod_3849 <- mkDebugOperation(mod_3849_inner, "mod_3849");
    Operation_IFC mod_3850_inner <- mkFlatten(0);
    Operation_IFC mod_3850 <- mkDebugOperation(mod_3850_inner, "mod_3850");
    Operation_IFC mod_3851_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3851 <- mkDebugOperation(mod_3851_inner, "mod_3851");
    Operation_IFC mod_3852_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3852 <- mkDebugOperation(mod_3852_inner, "mod_3852");
    PMU_IFC mod_3853_bufferize <- mkPMU(2);
    Operation_IFC mod_3853_inner = mod_3853_bufferize.operation;
    Operation_IFC mod_3853 <- mkDebugOperation(mod_3853_inner, "mod_3853");
    rule rule_4930;
        ChannelMessage t;
        t <- mod_3817.get(0);
        mod_3853.put(0, t);
    endrule
    rule rule_4931;
        ChannelMessage t;
        t <- mod_3841.get(0);
        mod_3842.put(0, t);
    endrule
    rule rule_4932;
        ChannelMessage t;
        t <- mod_3824.get(0);
        mod_3825.put(0, t);
    endrule
    rule rule_4933;
        ChannelMessage t;
        t <- mod_3852.get(0);
        mod_3819.put(1, t);
    endrule
    rule rule_4934;
        ChannelMessage t;
        t <- mod_3832.get(1);
        mod_3828.put(1, t);
    endrule
    rule rule_4935;
        ChannelMessage t;
        t <- mod_3853.get(1);
        mod_3817.put(1, t);
    endrule
    rule rule_4936;
        ChannelMessage t;
        t <- mod_3821.get(0);
        mod_3851.put(0, t);
    endrule
    rule rule_4937;
        ChannelMessage t;
        t <- mod_3816.get(0);
        mod_3817.put(0, t);
    endrule
    rule rule_4938;
        ChannelMessage t;
        t <- mod_3848.get(0);
        mod_3847.put(1, t);
    endrule
    rule rule_4939;
        ChannelMessage t;
        t <- mod_3818.get(3);
        mod_3819.put(0, t);
    endrule
    rule rule_4940;
        ChannelMessage t;
        t <- mod_3831.get(0);
        mod_3831.put(1, t);
    endrule
    rule rule_4941;
        ChannelMessage t;
        t <- mod_3831.get(1);
        mod_3829.put(1, t);
    endrule
    rule rule_4942;
        ChannelMessage t;
        t <- mod_3844.get(0);
        mod_3843.put(0, t);
    endrule
    rule rule_4943;
        ChannelMessage t;
        t <- mod_3819.get(0);
        mod_3852.put(0, t);
    endrule
    rule rule_4944;
        ChannelMessage t;
        t <- mod_3828.get(0);
        mod_3832.put(0, t);
    endrule
    rule rule_4945;
        ChannelMessage t;
        t <- mod_3825.get(1);
        mod_3826.put(0, t);
    endrule
    rule rule_4946;
        ChannelMessage t;
        t <- mod_3828.get(1);
        mod_3829.put(0, t);
    endrule
    rule rule_4947;
        ChannelMessage t;
        t <- mod_3840.get(0);
        mod_3839.put(0, t);
    endrule
    rule rule_4948;
        ChannelMessage t;
        t <- mod_3829.get(0);
        mod_3831.put(0, t);
    endrule
    rule rule_4949;
        ChannelMessage t;
        t <- mod_3820.get(0);
        mod_3845.put(0, t);
    endrule
    rule rule_4950;
        ChannelMessage t;
        t <- mod_3850.get(0);
        mod_3849.put(0, t);
    endrule
    rule rule_4951;
        ChannelMessage t;
        t <- mod_3833.get(1);
        mod_3826.put(1, t);
    endrule
    rule rule_4952;
        ChannelMessage t;
        t <- mod_3851.get(0);
        mod_3821.put(1, t);
    endrule
    rule rule_4953;
        ChannelMessage t;
        t <- mod_3847.get(1);
        mod_3822.put(1, t);
    endrule
    rule rule_4954;
        ChannelMessage t;
        t <- mod_3835.get(0);
        mod_3833.put(0, t);
    endrule
    rule rule_4955;
        ChannelMessage t;
        t <- mod_3819.get(1);
        mod_3820.put(0, t);
    endrule
    rule rule_4956;
        ChannelMessage t;
        t <- mod_3836.get(0);
        mod_3835.put(0, t);
    endrule
    rule rule_4957;
        ChannelMessage t;
        t <- mod_3846.get(0);
        mod_3845.put(1, t);
    endrule
    rule rule_4958;
        ChannelMessage t;
        t <- mod_3845.get(0);
        mod_3846.put(0, t);
    endrule
    rule rule_4959;
        ChannelMessage t;
        t <- mod_3823.get(0);
        mod_3824.put(0, t);
    endrule
    rule rule_4960;
        ChannelMessage t;
        t <- mod_3829.get(1);
        mod_3830.put(1, t);
    endrule
    rule rule_4961;
        ChannelMessage t;
        t <- mod_3839.get(0);
        mod_3838.put(0, t);
    endrule
    rule rule_4962;
        ChannelMessage t;
        t <- mod_3832.get(0);
        mod_3832.put(1, t);
    endrule
    rule rule_4963;
        ChannelMessage t;
        t <- mod_3843.get(0);
        mod_3841.put(0, t);
    endrule
    rule rule_4964;
        ChannelMessage t;
        t <- mod_3826.get(0);
        mod_3827.put(0, t);
    endrule
    rule rule_4965;
        ChannelMessage t;
        t <- mod_3853.get(0);
        mod_3853.put(1, t);
    endrule
    rule rule_4966;
        ChannelMessage t;
        t <- mod_3825.get(0);
        mod_3837.put(0, t);
    endrule
    rule rule_4967;
        ChannelMessage t;
        t <- mod_3842.get(0);
        mod_3841.put(1, t);
    endrule
    rule rule_4968;
        ChannelMessage t;
        t <- mod_3845.get(1);
        mod_3840.put(0, t);
    endrule
    rule rule_4969;
        ChannelMessage t;
        t <- mod_3847.get(0);
        mod_3848.put(0, t);
    endrule
    rule rule_4970;
        ChannelMessage t;
        t <- mod_3821.get(1);
        mod_3822.put(0, t);
    endrule
    rule rule_4971;
        ChannelMessage t;
        t <- mod_3834.get(0);
        mod_3833.put(1, t);
    endrule
    rule rule_4972;
        ChannelMessage t;
        t <- mod_3841.get(1);
        mod_3840.put(1, t);
    endrule
    rule rule_4973;
        ChannelMessage t;
        t <- mod_3815.get(0);
        mod_3816.put(0, t);
    endrule
    rule rule_4974;
        ChannelMessage t;
        t <- mod_3822.get(0);
        mod_3823.put(0, t);
    endrule
    rule rule_4975;
        ChannelMessage t;
        t <- mod_3817.get(1);
        mod_3818.put(0, t);
    endrule
    rule rule_4976;
        ChannelMessage t;
        t <- mod_3833.get(0);
        mod_3834.put(0, t);
    endrule
    rule rule_4977;
        ChannelMessage t;
        t <- mod_3849.get(0);
        mod_3847.put(0, t);
    endrule
    rule rule_4978;
        ChannelMessage t;
        t <- mod_3820.get(1);
        mod_3821.put(0, t);
    endrule
    rule rule_4979;
        ChannelMessage t;
        t <- mod_3814.get(0);
        mod_3815.put(0, t);
    endrule
    rule rule_4980;
        ChannelMessage t;
        t <- mod_3837.get(0);
        mod_3825.put(1, t);
    endrule
    rule rule_4981;
        ChannelMessage t;
        t <- mod_3838.get(0);
        mod_3824.put(1, t);
    endrule
    rule rule_4982;
        ChannelMessage t;
        t <- mod_3827.get(0);
        mod_3828.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3814.put(0, t);
        end
        if (i == 1) begin
            mod_3830.put(0, t);
        end
        if (i == 2) begin
            mod_3836.put(0, t);
        end
        if (i == 3) begin
            mod_3844.put(0, t);
        end
        if (i == 4) begin
            mod_3850.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 2) begin
            t <- mod_3818.get(0);
        end
        if (i == 1) begin
            t <- mod_3818.get(1);
        end
        if (i == 3) begin
            t <- mod_3818.get(2);
        end
        if (i == 0) begin
            t <- mod_3830.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6128 (Operation_IFC);
    Operation_IFC mod_3855_inner <- mkReshape(2, 64);
    Operation_IFC mod_3855 <- mkDebugOperation(mod_3855_inner, "mod_3855");
    Operation_IFC mod_3856_inner <- mkFlatten(1);
    Operation_IFC mod_3856 <- mkDebugOperation(mod_3856_inner, "mod_3856");
    Operation_IFC mod_3857_inner <- mkFlatten(2);
    Operation_IFC mod_3857 <- mkDebugOperation(mod_3857_inner, "mod_3857");
    Operation_IFC mod_3858_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3858 <- mkDebugOperation(mod_3858_inner, "mod_3858");
    Broadcast_IFC#(4) mod_3859_inner <- mkBroadcast(4);
    Operation_IFC mod_3859 <- mkDebugOperation(mod_3859_inner.op, "mod_3859");
    PMU_IFC mod_3860_bufferize <- mkPMU(2);
    Operation_IFC mod_3860_inner = mod_3860_bufferize.operation;
    Operation_IFC mod_3860 <- mkDebugOperation(mod_3860_inner, "mod_3860");
    Broadcast_IFC#(2) mod_3861_inner <- mkBroadcast(2);
    Operation_IFC mod_3861 <- mkDebugOperation(mod_3861_inner.op, "mod_3861");
    PMU_IFC mod_3862_bufferize <- mkPMU(1);
    Operation_IFC mod_3862_inner = mod_3862_bufferize.operation;
    Operation_IFC mod_3862 <- mkDebugOperation(mod_3862_inner, "mod_3862");
    Operation_IFC mod_3863_inner <- mkBinaryMap(1062, matmul_t_tile);
    Operation_IFC mod_3863 <- mkDebugOperation(mod_3863_inner, "mod_3863");
    Operation_IFC mod_3864_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3864 <- mkDebugOperation(mod_3864_inner, "mod_3864");
    Operation_IFC mod_3865_inner <- mkBinaryMap(1830, mul_tile);
    Operation_IFC mod_3865 <- mkDebugOperation(mod_3865_inner, "mod_3865");
    PMU_IFC mod_3866_bufferize <- mkPMU(1);
    Operation_IFC mod_3866_inner = mod_3866_bufferize.operation;
    Operation_IFC mod_3866 <- mkDebugOperation(mod_3866_inner, "mod_3866");
    Operation_IFC mod_3867_inner <- mkBinaryMap(2375, matmul_t_tile);
    Operation_IFC mod_3867 <- mkDebugOperation(mod_3867_inner, "mod_3867");
    Operation_IFC mod_3868_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3868 <- mkDebugOperation(mod_3868_inner, "mod_3868");
    Operation_IFC mod_3869_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3869 <- mkDebugOperation(mod_3869_inner, "mod_3869");
    Operation_IFC mod_3870_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3870 <- mkDebugOperation(mod_3870_inner, "mod_3870");
    Operation_IFC mod_3871_inner <- mkBinaryMap(2729, mul_tile);
    Operation_IFC mod_3871 <- mkDebugOperation(mod_3871_inner, "mod_3871");
    PMU_IFC mod_3872_bufferize <- mkPMU(1);
    Operation_IFC mod_3872_inner = mod_3872_bufferize.operation;
    Operation_IFC mod_3872 <- mkDebugOperation(mod_3872_inner, "mod_3872");
    PMU_IFC mod_3873_bufferize <- mkPMU(2);
    Operation_IFC mod_3873_inner = mod_3873_bufferize.operation;
    Operation_IFC mod_3873 <- mkDebugOperation(mod_3873_inner, "mod_3873");
    PMU_IFC mod_3874_bufferize <- mkPMU(2);
    Operation_IFC mod_3874_inner = mod_3874_bufferize.operation;
    Operation_IFC mod_3874 <- mkDebugOperation(mod_3874_inner, "mod_3874");
    Operation_IFC mod_3875_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3875 <- mkDebugOperation(mod_3875_inner, "mod_3875");
    Operation_IFC mod_3876_inner <- mkFlatten(1);
    Operation_IFC mod_3876 <- mkDebugOperation(mod_3876_inner, "mod_3876");
    Operation_IFC mod_3877_inner <- mkFlatten(0);
    Operation_IFC mod_3877 <- mkDebugOperation(mod_3877_inner, "mod_3877");
    Operation_IFC mod_3878_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3878 <- mkDebugOperation(mod_3878_inner, "mod_3878");
    Operation_IFC mod_3879_inner <- mkUnaryMap(1702, silu_tile);
    Operation_IFC mod_3879 <- mkDebugOperation(mod_3879_inner, "mod_3879");
    Operation_IFC mod_3880_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3880 <- mkDebugOperation(mod_3880_inner, "mod_3880");
    Operation_IFC mod_3881_inner <- mkBinaryMap(1574, matmul_t_tile);
    Operation_IFC mod_3881 <- mkDebugOperation(mod_3881_inner, "mod_3881");
    PMU_IFC mod_3882_bufferize <- mkPMU(2);
    Operation_IFC mod_3882_inner = mod_3882_bufferize.operation;
    Operation_IFC mod_3882 <- mkDebugOperation(mod_3882_inner, "mod_3882");
    Operation_IFC mod_3883_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3883 <- mkDebugOperation(mod_3883_inner, "mod_3883");
    Operation_IFC mod_3884_inner <- mkFlatten(1);
    Operation_IFC mod_3884 <- mkDebugOperation(mod_3884_inner, "mod_3884");
    Operation_IFC mod_3885_inner <- mkFlatten(0);
    Operation_IFC mod_3885 <- mkDebugOperation(mod_3885_inner, "mod_3885");
    PMU_IFC mod_3886_bufferize <- mkPMU(1);
    Operation_IFC mod_3886_inner = mod_3886_bufferize.operation;
    Operation_IFC mod_3886 <- mkDebugOperation(mod_3886_inner, "mod_3886");
    Operation_IFC mod_3887_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3887 <- mkDebugOperation(mod_3887_inner, "mod_3887");
    PMU_IFC mod_3888_bufferize <- mkPMU(2);
    Operation_IFC mod_3888_inner = mod_3888_bufferize.operation;
    Operation_IFC mod_3888 <- mkDebugOperation(mod_3888_inner, "mod_3888");
    Operation_IFC mod_3889_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3889 <- mkDebugOperation(mod_3889_inner, "mod_3889");
    Operation_IFC mod_3890_inner <- mkFlatten(1);
    Operation_IFC mod_3890 <- mkDebugOperation(mod_3890_inner, "mod_3890");
    Operation_IFC mod_3891_inner <- mkFlatten(0);
    Operation_IFC mod_3891 <- mkDebugOperation(mod_3891_inner, "mod_3891");
    Operation_IFC mod_3892_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3892 <- mkDebugOperation(mod_3892_inner, "mod_3892");
    Operation_IFC mod_3893_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3893 <- mkDebugOperation(mod_3893_inner, "mod_3893");
    PMU_IFC mod_3894_bufferize <- mkPMU(2);
    Operation_IFC mod_3894_inner = mod_3894_bufferize.operation;
    Operation_IFC mod_3894 <- mkDebugOperation(mod_3894_inner, "mod_3894");
    rule rule_4983;
        ChannelMessage t;
        t <- mod_3858.get(0);
        mod_3894.put(0, t);
    endrule
    rule rule_4984;
        ChannelMessage t;
        t <- mod_3883.get(0);
        mod_3882.put(1, t);
    endrule
    rule rule_4985;
        ChannelMessage t;
        t <- mod_3888.get(1);
        mod_3863.put(1, t);
    endrule
    rule rule_4986;
        ChannelMessage t;
        t <- mod_3869.get(1);
        mod_3870.put(0, t);
    endrule
    rule rule_4987;
        ChannelMessage t;
        t <- mod_3882.get(0);
        mod_3883.put(0, t);
    endrule
    rule rule_4988;
        ChannelMessage t;
        t <- mod_3855.get(0);
        mod_3856.put(0, t);
    endrule
    rule rule_4989;
        ChannelMessage t;
        t <- mod_3869.get(0);
        mod_3873.put(0, t);
    endrule
    rule rule_4990;
        ChannelMessage t;
        t <- mod_3863.get(0);
        mod_3864.put(0, t);
    endrule
    rule rule_4991;
        ChannelMessage t;
        t <- mod_3890.get(0);
        mod_3888.put(0, t);
    endrule
    rule rule_4992;
        ChannelMessage t;
        t <- mod_3878.get(0);
        mod_3866.put(1, t);
    endrule
    rule rule_4993;
        ChannelMessage t;
        t <- mod_3886.get(1);
        mod_3881.put(0, t);
    endrule
    rule rule_4994;
        ChannelMessage t;
        t <- mod_3870.get(1);
        mod_3871.put(1, t);
    endrule
    rule rule_4995;
        ChannelMessage t;
        t <- mod_3860.get(0);
        mod_3893.put(0, t);
    endrule
    rule rule_4996;
        ChannelMessage t;
        t <- mod_3859.get(3);
        mod_3860.put(0, t);
    endrule
    rule rule_4997;
        ChannelMessage t;
        t <- mod_3885.get(0);
        mod_3884.put(0, t);
    endrule
    rule rule_4998;
        ChannelMessage t;
        t <- mod_3861.get(1);
        mod_3862.put(0, t);
    endrule
    rule rule_4999;
        ChannelMessage t;
        t <- mod_3873.get(1);
        mod_3869.put(1, t);
    endrule
    rule rule_5000;
        ChannelMessage t;
        t <- mod_3880.get(0);
        mod_3879.put(0, t);
    endrule
    rule rule_5001;
        ChannelMessage t;
        t <- mod_3866.get(1);
        mod_3867.put(0, t);
    endrule
    rule rule_5002;
        ChannelMessage t;
        t <- mod_3881.get(0);
        mod_3880.put(0, t);
    endrule
    rule rule_5003;
        ChannelMessage t;
        t <- mod_3882.get(1);
        mod_3881.put(1, t);
    endrule
    rule rule_5004;
        ChannelMessage t;
        t <- mod_3857.get(0);
        mod_3858.put(0, t);
    endrule
    rule rule_5005;
        ChannelMessage t;
        t <- mod_3894.get(1);
        mod_3858.put(1, t);
    endrule
    rule rule_5006;
        ChannelMessage t;
        t <- mod_3870.get(0);
        mod_3872.put(0, t);
    endrule
    rule rule_5007;
        ChannelMessage t;
        t <- mod_3862.get(0);
        mod_3892.put(0, t);
    endrule
    rule rule_5008;
        ChannelMessage t;
        t <- mod_3876.get(0);
        mod_3874.put(0, t);
    endrule
    rule rule_5009;
        ChannelMessage t;
        t <- mod_3884.get(0);
        mod_3882.put(0, t);
    endrule
    rule rule_5010;
        ChannelMessage t;
        t <- mod_3860.get(1);
        mod_3861.put(0, t);
    endrule
    rule rule_5011;
        ChannelMessage t;
        t <- mod_3862.get(1);
        mod_3863.put(0, t);
    endrule
    rule rule_5012;
        ChannelMessage t;
        t <- mod_3872.get(0);
        mod_3872.put(1, t);
    endrule
    rule rule_5013;
        ChannelMessage t;
        t <- mod_3879.get(0);
        mod_3865.put(1, t);
    endrule
    rule rule_5014;
        ChannelMessage t;
        t <- mod_3892.get(0);
        mod_3862.put(1, t);
    endrule
    rule rule_5015;
        ChannelMessage t;
        t <- mod_3893.get(0);
        mod_3860.put(1, t);
    endrule
    rule rule_5016;
        ChannelMessage t;
        t <- mod_3867.get(0);
        mod_3868.put(0, t);
    endrule
    rule rule_5017;
        ChannelMessage t;
        t <- mod_3891.get(0);
        mod_3890.put(0, t);
    endrule
    rule rule_5018;
        ChannelMessage t;
        t <- mod_3875.get(0);
        mod_3874.put(1, t);
    endrule
    rule rule_5019;
        ChannelMessage t;
        t <- mod_3873.get(0);
        mod_3873.put(1, t);
    endrule
    rule rule_5020;
        ChannelMessage t;
        t <- mod_3864.get(0);
        mod_3865.put(0, t);
    endrule
    rule rule_5021;
        ChannelMessage t;
        t <- mod_3865.get(0);
        mod_3866.put(0, t);
    endrule
    rule rule_5022;
        ChannelMessage t;
        t <- mod_3877.get(0);
        mod_3876.put(0, t);
    endrule
    rule rule_5023;
        ChannelMessage t;
        t <- mod_3858.get(1);
        mod_3859.put(0, t);
    endrule
    rule rule_5024;
        ChannelMessage t;
        t <- mod_3894.get(0);
        mod_3894.put(1, t);
    endrule
    rule rule_5025;
        ChannelMessage t;
        t <- mod_3886.get(0);
        mod_3887.put(0, t);
    endrule
    rule rule_5026;
        ChannelMessage t;
        t <- mod_3868.get(0);
        mod_3869.put(0, t);
    endrule
    rule rule_5027;
        ChannelMessage t;
        t <- mod_3889.get(0);
        mod_3888.put(1, t);
    endrule
    rule rule_5028;
        ChannelMessage t;
        t <- mod_3866.get(0);
        mod_3878.put(0, t);
    endrule
    rule rule_5029;
        ChannelMessage t;
        t <- mod_3888.get(0);
        mod_3889.put(0, t);
    endrule
    rule rule_5030;
        ChannelMessage t;
        t <- mod_3861.get(0);
        mod_3886.put(0, t);
    endrule
    rule rule_5031;
        ChannelMessage t;
        t <- mod_3856.get(0);
        mod_3857.put(0, t);
    endrule
    rule rule_5032;
        ChannelMessage t;
        t <- mod_3874.get(0);
        mod_3875.put(0, t);
    endrule
    rule rule_5033;
        ChannelMessage t;
        t <- mod_3887.get(0);
        mod_3886.put(1, t);
    endrule
    rule rule_5034;
        ChannelMessage t;
        t <- mod_3874.get(1);
        mod_3867.put(1, t);
    endrule
    rule rule_5035;
        ChannelMessage t;
        t <- mod_3872.get(1);
        mod_3870.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3855.put(0, t);
        end
        if (i == 1) begin
            mod_3871.put(0, t);
        end
        if (i == 2) begin
            mod_3877.put(0, t);
        end
        if (i == 3) begin
            mod_3885.put(0, t);
        end
        if (i == 4) begin
            mod_3891.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_3859.get(0);
        end
        if (i == 3) begin
            t <- mod_3859.get(1);
        end
        if (i == 1) begin
            t <- mod_3859.get(2);
        end
        if (i == 2) begin
            t <- mod_3871.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6129 (Operation_IFC);
    Operation_IFC mod_3896_inner <- mkReshape(2, 64);
    Operation_IFC mod_3896 <- mkDebugOperation(mod_3896_inner, "mod_3896");
    Operation_IFC mod_3897_inner <- mkFlatten(1);
    Operation_IFC mod_3897 <- mkDebugOperation(mod_3897_inner, "mod_3897");
    Operation_IFC mod_3898_inner <- mkFlatten(2);
    Operation_IFC mod_3898 <- mkDebugOperation(mod_3898_inner, "mod_3898");
    Operation_IFC mod_3899_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3899 <- mkDebugOperation(mod_3899_inner, "mod_3899");
    Broadcast_IFC#(4) mod_3900_inner <- mkBroadcast(4);
    Operation_IFC mod_3900 <- mkDebugOperation(mod_3900_inner.op, "mod_3900");
    PMU_IFC mod_3901_bufferize <- mkPMU(2);
    Operation_IFC mod_3901_inner = mod_3901_bufferize.operation;
    Operation_IFC mod_3901 <- mkDebugOperation(mod_3901_inner, "mod_3901");
    Broadcast_IFC#(2) mod_3902_inner <- mkBroadcast(2);
    Operation_IFC mod_3902 <- mkDebugOperation(mod_3902_inner.op, "mod_3902");
    PMU_IFC mod_3903_bufferize <- mkPMU(1);
    Operation_IFC mod_3903_inner = mod_3903_bufferize.operation;
    Operation_IFC mod_3903 <- mkDebugOperation(mod_3903_inner, "mod_3903");
    Operation_IFC mod_3904_inner <- mkBinaryMap(1061, matmul_t_tile);
    Operation_IFC mod_3904 <- mkDebugOperation(mod_3904_inner, "mod_3904");
    Operation_IFC mod_3905_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3905 <- mkDebugOperation(mod_3905_inner, "mod_3905");
    Operation_IFC mod_3906_inner <- mkBinaryMap(1829, mul_tile);
    Operation_IFC mod_3906 <- mkDebugOperation(mod_3906_inner, "mod_3906");
    PMU_IFC mod_3907_bufferize <- mkPMU(1);
    Operation_IFC mod_3907_inner = mod_3907_bufferize.operation;
    Operation_IFC mod_3907 <- mkDebugOperation(mod_3907_inner, "mod_3907");
    Operation_IFC mod_3908_inner <- mkBinaryMap(2373, matmul_t_tile);
    Operation_IFC mod_3908 <- mkDebugOperation(mod_3908_inner, "mod_3908");
    Operation_IFC mod_3909_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3909 <- mkDebugOperation(mod_3909_inner, "mod_3909");
    Operation_IFC mod_3910_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3910 <- mkDebugOperation(mod_3910_inner, "mod_3910");
    Operation_IFC mod_3911_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3911 <- mkDebugOperation(mod_3911_inner, "mod_3911");
    Operation_IFC mod_3912_inner <- mkBinaryMap(2728, mul_tile);
    Operation_IFC mod_3912 <- mkDebugOperation(mod_3912_inner, "mod_3912");
    PMU_IFC mod_3913_bufferize <- mkPMU(1);
    Operation_IFC mod_3913_inner = mod_3913_bufferize.operation;
    Operation_IFC mod_3913 <- mkDebugOperation(mod_3913_inner, "mod_3913");
    PMU_IFC mod_3914_bufferize <- mkPMU(2);
    Operation_IFC mod_3914_inner = mod_3914_bufferize.operation;
    Operation_IFC mod_3914 <- mkDebugOperation(mod_3914_inner, "mod_3914");
    PMU_IFC mod_3915_bufferize <- mkPMU(2);
    Operation_IFC mod_3915_inner = mod_3915_bufferize.operation;
    Operation_IFC mod_3915 <- mkDebugOperation(mod_3915_inner, "mod_3915");
    Operation_IFC mod_3916_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3916 <- mkDebugOperation(mod_3916_inner, "mod_3916");
    Operation_IFC mod_3917_inner <- mkFlatten(1);
    Operation_IFC mod_3917 <- mkDebugOperation(mod_3917_inner, "mod_3917");
    Operation_IFC mod_3918_inner <- mkFlatten(0);
    Operation_IFC mod_3918 <- mkDebugOperation(mod_3918_inner, "mod_3918");
    Operation_IFC mod_3919_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3919 <- mkDebugOperation(mod_3919_inner, "mod_3919");
    Operation_IFC mod_3920_inner <- mkUnaryMap(1701, silu_tile);
    Operation_IFC mod_3920 <- mkDebugOperation(mod_3920_inner, "mod_3920");
    Operation_IFC mod_3921_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3921 <- mkDebugOperation(mod_3921_inner, "mod_3921");
    Operation_IFC mod_3922_inner <- mkBinaryMap(1573, matmul_t_tile);
    Operation_IFC mod_3922 <- mkDebugOperation(mod_3922_inner, "mod_3922");
    PMU_IFC mod_3923_bufferize <- mkPMU(2);
    Operation_IFC mod_3923_inner = mod_3923_bufferize.operation;
    Operation_IFC mod_3923 <- mkDebugOperation(mod_3923_inner, "mod_3923");
    Operation_IFC mod_3924_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3924 <- mkDebugOperation(mod_3924_inner, "mod_3924");
    Operation_IFC mod_3925_inner <- mkFlatten(1);
    Operation_IFC mod_3925 <- mkDebugOperation(mod_3925_inner, "mod_3925");
    Operation_IFC mod_3926_inner <- mkFlatten(0);
    Operation_IFC mod_3926 <- mkDebugOperation(mod_3926_inner, "mod_3926");
    PMU_IFC mod_3927_bufferize <- mkPMU(1);
    Operation_IFC mod_3927_inner = mod_3927_bufferize.operation;
    Operation_IFC mod_3927 <- mkDebugOperation(mod_3927_inner, "mod_3927");
    Operation_IFC mod_3928_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3928 <- mkDebugOperation(mod_3928_inner, "mod_3928");
    PMU_IFC mod_3929_bufferize <- mkPMU(2);
    Operation_IFC mod_3929_inner = mod_3929_bufferize.operation;
    Operation_IFC mod_3929 <- mkDebugOperation(mod_3929_inner, "mod_3929");
    Operation_IFC mod_3930_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3930 <- mkDebugOperation(mod_3930_inner, "mod_3930");
    Operation_IFC mod_3931_inner <- mkFlatten(1);
    Operation_IFC mod_3931 <- mkDebugOperation(mod_3931_inner, "mod_3931");
    Operation_IFC mod_3932_inner <- mkFlatten(0);
    Operation_IFC mod_3932 <- mkDebugOperation(mod_3932_inner, "mod_3932");
    Operation_IFC mod_3933_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3933 <- mkDebugOperation(mod_3933_inner, "mod_3933");
    Operation_IFC mod_3934_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3934 <- mkDebugOperation(mod_3934_inner, "mod_3934");
    PMU_IFC mod_3935_bufferize <- mkPMU(2);
    Operation_IFC mod_3935_inner = mod_3935_bufferize.operation;
    Operation_IFC mod_3935 <- mkDebugOperation(mod_3935_inner, "mod_3935");
    rule rule_5036;
        ChannelMessage t;
        t <- mod_3920.get(0);
        mod_3906.put(1, t);
    endrule
    rule rule_5037;
        ChannelMessage t;
        t <- mod_3924.get(0);
        mod_3923.put(1, t);
    endrule
    rule rule_5038;
        ChannelMessage t;
        t <- mod_3917.get(0);
        mod_3915.put(0, t);
    endrule
    rule rule_5039;
        ChannelMessage t;
        t <- mod_3927.get(0);
        mod_3928.put(0, t);
    endrule
    rule rule_5040;
        ChannelMessage t;
        t <- mod_3896.get(0);
        mod_3897.put(0, t);
    endrule
    rule rule_5041;
        ChannelMessage t;
        t <- mod_3930.get(0);
        mod_3929.put(1, t);
    endrule
    rule rule_5042;
        ChannelMessage t;
        t <- mod_3921.get(0);
        mod_3920.put(0, t);
    endrule
    rule rule_5043;
        ChannelMessage t;
        t <- mod_3918.get(0);
        mod_3917.put(0, t);
    endrule
    rule rule_5044;
        ChannelMessage t;
        t <- mod_3897.get(0);
        mod_3898.put(0, t);
    endrule
    rule rule_5045;
        ChannelMessage t;
        t <- mod_3929.get(1);
        mod_3904.put(1, t);
    endrule
    rule rule_5046;
        ChannelMessage t;
        t <- mod_3904.get(0);
        mod_3905.put(0, t);
    endrule
    rule rule_5047;
        ChannelMessage t;
        t <- mod_3911.get(1);
        mod_3912.put(1, t);
    endrule
    rule rule_5048;
        ChannelMessage t;
        t <- mod_3910.get(0);
        mod_3914.put(0, t);
    endrule
    rule rule_5049;
        ChannelMessage t;
        t <- mod_3907.get(0);
        mod_3919.put(0, t);
    endrule
    rule rule_5050;
        ChannelMessage t;
        t <- mod_3914.get(1);
        mod_3910.put(1, t);
    endrule
    rule rule_5051;
        ChannelMessage t;
        t <- mod_3909.get(0);
        mod_3910.put(0, t);
    endrule
    rule rule_5052;
        ChannelMessage t;
        t <- mod_3913.get(1);
        mod_3911.put(1, t);
    endrule
    rule rule_5053;
        ChannelMessage t;
        t <- mod_3908.get(0);
        mod_3909.put(0, t);
    endrule
    rule rule_5054;
        ChannelMessage t;
        t <- mod_3929.get(0);
        mod_3930.put(0, t);
    endrule
    rule rule_5055;
        ChannelMessage t;
        t <- mod_3899.get(0);
        mod_3935.put(0, t);
    endrule
    rule rule_5056;
        ChannelMessage t;
        t <- mod_3928.get(0);
        mod_3927.put(1, t);
    endrule
    rule rule_5057;
        ChannelMessage t;
        t <- mod_3914.get(0);
        mod_3914.put(1, t);
    endrule
    rule rule_5058;
        ChannelMessage t;
        t <- mod_3907.get(1);
        mod_3908.put(0, t);
    endrule
    rule rule_5059;
        ChannelMessage t;
        t <- mod_3903.get(1);
        mod_3904.put(0, t);
    endrule
    rule rule_5060;
        ChannelMessage t;
        t <- mod_3933.get(0);
        mod_3903.put(1, t);
    endrule
    rule rule_5061;
        ChannelMessage t;
        t <- mod_3901.get(1);
        mod_3902.put(0, t);
    endrule
    rule rule_5062;
        ChannelMessage t;
        t <- mod_3923.get(0);
        mod_3924.put(0, t);
    endrule
    rule rule_5063;
        ChannelMessage t;
        t <- mod_3910.get(1);
        mod_3911.put(0, t);
    endrule
    rule rule_5064;
        ChannelMessage t;
        t <- mod_3911.get(0);
        mod_3913.put(0, t);
    endrule
    rule rule_5065;
        ChannelMessage t;
        t <- mod_3902.get(0);
        mod_3927.put(0, t);
    endrule
    rule rule_5066;
        ChannelMessage t;
        t <- mod_3923.get(1);
        mod_3922.put(1, t);
    endrule
    rule rule_5067;
        ChannelMessage t;
        t <- mod_3925.get(0);
        mod_3923.put(0, t);
    endrule
    rule rule_5068;
        ChannelMessage t;
        t <- mod_3916.get(0);
        mod_3915.put(1, t);
    endrule
    rule rule_5069;
        ChannelMessage t;
        t <- mod_3905.get(0);
        mod_3906.put(0, t);
    endrule
    rule rule_5070;
        ChannelMessage t;
        t <- mod_3932.get(0);
        mod_3931.put(0, t);
    endrule
    rule rule_5071;
        ChannelMessage t;
        t <- mod_3931.get(0);
        mod_3929.put(0, t);
    endrule
    rule rule_5072;
        ChannelMessage t;
        t <- mod_3915.get(1);
        mod_3908.put(1, t);
    endrule
    rule rule_5073;
        ChannelMessage t;
        t <- mod_3913.get(0);
        mod_3913.put(1, t);
    endrule
    rule rule_5074;
        ChannelMessage t;
        t <- mod_3915.get(0);
        mod_3916.put(0, t);
    endrule
    rule rule_5075;
        ChannelMessage t;
        t <- mod_3901.get(0);
        mod_3934.put(0, t);
    endrule
    rule rule_5076;
        ChannelMessage t;
        t <- mod_3906.get(0);
        mod_3907.put(0, t);
    endrule
    rule rule_5077;
        ChannelMessage t;
        t <- mod_3900.get(3);
        mod_3901.put(0, t);
    endrule
    rule rule_5078;
        ChannelMessage t;
        t <- mod_3902.get(1);
        mod_3903.put(0, t);
    endrule
    rule rule_5079;
        ChannelMessage t;
        t <- mod_3903.get(0);
        mod_3933.put(0, t);
    endrule
    rule rule_5080;
        ChannelMessage t;
        t <- mod_3898.get(0);
        mod_3899.put(0, t);
    endrule
    rule rule_5081;
        ChannelMessage t;
        t <- mod_3927.get(1);
        mod_3922.put(0, t);
    endrule
    rule rule_5082;
        ChannelMessage t;
        t <- mod_3926.get(0);
        mod_3925.put(0, t);
    endrule
    rule rule_5083;
        ChannelMessage t;
        t <- mod_3934.get(0);
        mod_3901.put(1, t);
    endrule
    rule rule_5084;
        ChannelMessage t;
        t <- mod_3935.get(1);
        mod_3899.put(1, t);
    endrule
    rule rule_5085;
        ChannelMessage t;
        t <- mod_3922.get(0);
        mod_3921.put(0, t);
    endrule
    rule rule_5086;
        ChannelMessage t;
        t <- mod_3899.get(1);
        mod_3900.put(0, t);
    endrule
    rule rule_5087;
        ChannelMessage t;
        t <- mod_3919.get(0);
        mod_3907.put(1, t);
    endrule
    rule rule_5088;
        ChannelMessage t;
        t <- mod_3935.get(0);
        mod_3935.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3896.put(0, t);
        end
        if (i == 1) begin
            mod_3912.put(0, t);
        end
        if (i == 2) begin
            mod_3918.put(0, t);
        end
        if (i == 3) begin
            mod_3926.put(0, t);
        end
        if (i == 4) begin
            mod_3932.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_3900.get(0);
        end
        if (i == 3) begin
            t <- mod_3900.get(1);
        end
        if (i == 2) begin
            t <- mod_3900.get(2);
        end
        if (i == 0) begin
            t <- mod_3912.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6130 (Operation_IFC);
    Operation_IFC mod_3937_inner <- mkReshape(2, 64);
    Operation_IFC mod_3937 <- mkDebugOperation(mod_3937_inner, "mod_3937");
    Operation_IFC mod_3938_inner <- mkFlatten(1);
    Operation_IFC mod_3938 <- mkDebugOperation(mod_3938_inner, "mod_3938");
    Operation_IFC mod_3939_inner <- mkFlatten(2);
    Operation_IFC mod_3939 <- mkDebugOperation(mod_3939_inner, "mod_3939");
    Operation_IFC mod_3940_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3940 <- mkDebugOperation(mod_3940_inner, "mod_3940");
    Broadcast_IFC#(4) mod_3941_inner <- mkBroadcast(4);
    Operation_IFC mod_3941 <- mkDebugOperation(mod_3941_inner.op, "mod_3941");
    PMU_IFC mod_3942_bufferize <- mkPMU(2);
    Operation_IFC mod_3942_inner = mod_3942_bufferize.operation;
    Operation_IFC mod_3942 <- mkDebugOperation(mod_3942_inner, "mod_3942");
    Broadcast_IFC#(2) mod_3943_inner <- mkBroadcast(2);
    Operation_IFC mod_3943 <- mkDebugOperation(mod_3943_inner.op, "mod_3943");
    PMU_IFC mod_3944_bufferize <- mkPMU(1);
    Operation_IFC mod_3944_inner = mod_3944_bufferize.operation;
    Operation_IFC mod_3944 <- mkDebugOperation(mod_3944_inner, "mod_3944");
    Operation_IFC mod_3945_inner <- mkBinaryMap(1060, matmul_t_tile);
    Operation_IFC mod_3945 <- mkDebugOperation(mod_3945_inner, "mod_3945");
    Operation_IFC mod_3946_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3946 <- mkDebugOperation(mod_3946_inner, "mod_3946");
    Operation_IFC mod_3947_inner <- mkBinaryMap(1828, mul_tile);
    Operation_IFC mod_3947 <- mkDebugOperation(mod_3947_inner, "mod_3947");
    PMU_IFC mod_3948_bufferize <- mkPMU(1);
    Operation_IFC mod_3948_inner = mod_3948_bufferize.operation;
    Operation_IFC mod_3948 <- mkDebugOperation(mod_3948_inner, "mod_3948");
    Operation_IFC mod_3949_inner <- mkBinaryMap(2371, matmul_t_tile);
    Operation_IFC mod_3949 <- mkDebugOperation(mod_3949_inner, "mod_3949");
    Operation_IFC mod_3950_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3950 <- mkDebugOperation(mod_3950_inner, "mod_3950");
    Operation_IFC mod_3951_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3951 <- mkDebugOperation(mod_3951_inner, "mod_3951");
    Operation_IFC mod_3952_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3952 <- mkDebugOperation(mod_3952_inner, "mod_3952");
    Operation_IFC mod_3953_inner <- mkBinaryMap(2727, mul_tile);
    Operation_IFC mod_3953 <- mkDebugOperation(mod_3953_inner, "mod_3953");
    PMU_IFC mod_3954_bufferize <- mkPMU(1);
    Operation_IFC mod_3954_inner = mod_3954_bufferize.operation;
    Operation_IFC mod_3954 <- mkDebugOperation(mod_3954_inner, "mod_3954");
    PMU_IFC mod_3955_bufferize <- mkPMU(2);
    Operation_IFC mod_3955_inner = mod_3955_bufferize.operation;
    Operation_IFC mod_3955 <- mkDebugOperation(mod_3955_inner, "mod_3955");
    PMU_IFC mod_3956_bufferize <- mkPMU(2);
    Operation_IFC mod_3956_inner = mod_3956_bufferize.operation;
    Operation_IFC mod_3956 <- mkDebugOperation(mod_3956_inner, "mod_3956");
    Operation_IFC mod_3957_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3957 <- mkDebugOperation(mod_3957_inner, "mod_3957");
    Operation_IFC mod_3958_inner <- mkFlatten(1);
    Operation_IFC mod_3958 <- mkDebugOperation(mod_3958_inner, "mod_3958");
    Operation_IFC mod_3959_inner <- mkFlatten(0);
    Operation_IFC mod_3959 <- mkDebugOperation(mod_3959_inner, "mod_3959");
    Operation_IFC mod_3960_inner <- mkRepeatStatic(3);
    Operation_IFC mod_3960 <- mkDebugOperation(mod_3960_inner, "mod_3960");
    Operation_IFC mod_3961_inner <- mkUnaryMap(1700, silu_tile);
    Operation_IFC mod_3961 <- mkDebugOperation(mod_3961_inner, "mod_3961");
    Operation_IFC mod_3962_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3962 <- mkDebugOperation(mod_3962_inner, "mod_3962");
    Operation_IFC mod_3963_inner <- mkBinaryMap(1572, matmul_t_tile);
    Operation_IFC mod_3963 <- mkDebugOperation(mod_3963_inner, "mod_3963");
    PMU_IFC mod_3964_bufferize <- mkPMU(2);
    Operation_IFC mod_3964_inner = mod_3964_bufferize.operation;
    Operation_IFC mod_3964 <- mkDebugOperation(mod_3964_inner, "mod_3964");
    Operation_IFC mod_3965_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3965 <- mkDebugOperation(mod_3965_inner, "mod_3965");
    Operation_IFC mod_3966_inner <- mkFlatten(1);
    Operation_IFC mod_3966 <- mkDebugOperation(mod_3966_inner, "mod_3966");
    Operation_IFC mod_3967_inner <- mkFlatten(0);
    Operation_IFC mod_3967 <- mkDebugOperation(mod_3967_inner, "mod_3967");
    PMU_IFC mod_3968_bufferize <- mkPMU(1);
    Operation_IFC mod_3968_inner = mod_3968_bufferize.operation;
    Operation_IFC mod_3968 <- mkDebugOperation(mod_3968_inner, "mod_3968");
    Operation_IFC mod_3969_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3969 <- mkDebugOperation(mod_3969_inner, "mod_3969");
    PMU_IFC mod_3970_bufferize <- mkPMU(2);
    Operation_IFC mod_3970_inner = mod_3970_bufferize.operation;
    Operation_IFC mod_3970 <- mkDebugOperation(mod_3970_inner, "mod_3970");
    Operation_IFC mod_3971_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3971 <- mkDebugOperation(mod_3971_inner, "mod_3971");
    Operation_IFC mod_3972_inner <- mkFlatten(1);
    Operation_IFC mod_3972 <- mkDebugOperation(mod_3972_inner, "mod_3972");
    Operation_IFC mod_3973_inner <- mkFlatten(0);
    Operation_IFC mod_3973 <- mkDebugOperation(mod_3973_inner, "mod_3973");
    Operation_IFC mod_3974_inner <- mkRepeatStatic(16);
    Operation_IFC mod_3974 <- mkDebugOperation(mod_3974_inner, "mod_3974");
    Operation_IFC mod_3975_inner <- mkRepeatStatic(2);
    Operation_IFC mod_3975 <- mkDebugOperation(mod_3975_inner, "mod_3975");
    PMU_IFC mod_3976_bufferize <- mkPMU(2);
    Operation_IFC mod_3976_inner = mod_3976_bufferize.operation;
    Operation_IFC mod_3976 <- mkDebugOperation(mod_3976_inner, "mod_3976");
    rule rule_5089;
        ChannelMessage t;
        t <- mod_3968.get(0);
        mod_3969.put(0, t);
    endrule
    rule rule_5090;
        ChannelMessage t;
        t <- mod_3951.get(1);
        mod_3952.put(0, t);
    endrule
    rule rule_5091;
        ChannelMessage t;
        t <- mod_3937.get(0);
        mod_3938.put(0, t);
    endrule
    rule rule_5092;
        ChannelMessage t;
        t <- mod_3944.get(0);
        mod_3974.put(0, t);
    endrule
    rule rule_5093;
        ChannelMessage t;
        t <- mod_3939.get(0);
        mod_3940.put(0, t);
    endrule
    rule rule_5094;
        ChannelMessage t;
        t <- mod_3972.get(0);
        mod_3970.put(0, t);
    endrule
    rule rule_5095;
        ChannelMessage t;
        t <- mod_3961.get(0);
        mod_3947.put(1, t);
    endrule
    rule rule_5096;
        ChannelMessage t;
        t <- mod_3956.get(1);
        mod_3949.put(1, t);
    endrule
    rule rule_5097;
        ChannelMessage t;
        t <- mod_3962.get(0);
        mod_3961.put(0, t);
    endrule
    rule rule_5098;
        ChannelMessage t;
        t <- mod_3964.get(0);
        mod_3965.put(0, t);
    endrule
    rule rule_5099;
        ChannelMessage t;
        t <- mod_3960.get(0);
        mod_3948.put(1, t);
    endrule
    rule rule_5100;
        ChannelMessage t;
        t <- mod_3950.get(0);
        mod_3951.put(0, t);
    endrule
    rule rule_5101;
        ChannelMessage t;
        t <- mod_3976.get(1);
        mod_3940.put(1, t);
    endrule
    rule rule_5102;
        ChannelMessage t;
        t <- mod_3940.get(0);
        mod_3976.put(0, t);
    endrule
    rule rule_5103;
        ChannelMessage t;
        t <- mod_3947.get(0);
        mod_3948.put(0, t);
    endrule
    rule rule_5104;
        ChannelMessage t;
        t <- mod_3957.get(0);
        mod_3956.put(1, t);
    endrule
    rule rule_5105;
        ChannelMessage t;
        t <- mod_3942.get(0);
        mod_3975.put(0, t);
    endrule
    rule rule_5106;
        ChannelMessage t;
        t <- mod_3943.get(1);
        mod_3944.put(0, t);
    endrule
    rule rule_5107;
        ChannelMessage t;
        t <- mod_3952.get(0);
        mod_3954.put(0, t);
    endrule
    rule rule_5108;
        ChannelMessage t;
        t <- mod_3971.get(0);
        mod_3970.put(1, t);
    endrule
    rule rule_5109;
        ChannelMessage t;
        t <- mod_3954.get(1);
        mod_3952.put(1, t);
    endrule
    rule rule_5110;
        ChannelMessage t;
        t <- mod_3964.get(1);
        mod_3963.put(1, t);
    endrule
    rule rule_5111;
        ChannelMessage t;
        t <- mod_3943.get(0);
        mod_3968.put(0, t);
    endrule
    rule rule_5112;
        ChannelMessage t;
        t <- mod_3955.get(0);
        mod_3955.put(1, t);
    endrule
    rule rule_5113;
        ChannelMessage t;
        t <- mod_3952.get(1);
        mod_3953.put(1, t);
    endrule
    rule rule_5114;
        ChannelMessage t;
        t <- mod_3970.get(0);
        mod_3971.put(0, t);
    endrule
    rule rule_5115;
        ChannelMessage t;
        t <- mod_3974.get(0);
        mod_3944.put(1, t);
    endrule
    rule rule_5116;
        ChannelMessage t;
        t <- mod_3941.get(3);
        mod_3942.put(0, t);
    endrule
    rule rule_5117;
        ChannelMessage t;
        t <- mod_3948.get(0);
        mod_3960.put(0, t);
    endrule
    rule rule_5118;
        ChannelMessage t;
        t <- mod_3949.get(0);
        mod_3950.put(0, t);
    endrule
    rule rule_5119;
        ChannelMessage t;
        t <- mod_3958.get(0);
        mod_3956.put(0, t);
    endrule
    rule rule_5120;
        ChannelMessage t;
        t <- mod_3969.get(0);
        mod_3968.put(1, t);
    endrule
    rule rule_5121;
        ChannelMessage t;
        t <- mod_3975.get(0);
        mod_3942.put(1, t);
    endrule
    rule rule_5122;
        ChannelMessage t;
        t <- mod_3945.get(0);
        mod_3946.put(0, t);
    endrule
    rule rule_5123;
        ChannelMessage t;
        t <- mod_3967.get(0);
        mod_3966.put(0, t);
    endrule
    rule rule_5124;
        ChannelMessage t;
        t <- mod_3944.get(1);
        mod_3945.put(0, t);
    endrule
    rule rule_5125;
        ChannelMessage t;
        t <- mod_3965.get(0);
        mod_3964.put(1, t);
    endrule
    rule rule_5126;
        ChannelMessage t;
        t <- mod_3976.get(0);
        mod_3976.put(1, t);
    endrule
    rule rule_5127;
        ChannelMessage t;
        t <- mod_3968.get(1);
        mod_3963.put(0, t);
    endrule
    rule rule_5128;
        ChannelMessage t;
        t <- mod_3954.get(0);
        mod_3954.put(1, t);
    endrule
    rule rule_5129;
        ChannelMessage t;
        t <- mod_3973.get(0);
        mod_3972.put(0, t);
    endrule
    rule rule_5130;
        ChannelMessage t;
        t <- mod_3940.get(1);
        mod_3941.put(0, t);
    endrule
    rule rule_5131;
        ChannelMessage t;
        t <- mod_3966.get(0);
        mod_3964.put(0, t);
    endrule
    rule rule_5132;
        ChannelMessage t;
        t <- mod_3942.get(1);
        mod_3943.put(0, t);
    endrule
    rule rule_5133;
        ChannelMessage t;
        t <- mod_3946.get(0);
        mod_3947.put(0, t);
    endrule
    rule rule_5134;
        ChannelMessage t;
        t <- mod_3955.get(1);
        mod_3951.put(1, t);
    endrule
    rule rule_5135;
        ChannelMessage t;
        t <- mod_3948.get(1);
        mod_3949.put(0, t);
    endrule
    rule rule_5136;
        ChannelMessage t;
        t <- mod_3938.get(0);
        mod_3939.put(0, t);
    endrule
    rule rule_5137;
        ChannelMessage t;
        t <- mod_3963.get(0);
        mod_3962.put(0, t);
    endrule
    rule rule_5138;
        ChannelMessage t;
        t <- mod_3956.get(0);
        mod_3957.put(0, t);
    endrule
    rule rule_5139;
        ChannelMessage t;
        t <- mod_3959.get(0);
        mod_3958.put(0, t);
    endrule
    rule rule_5140;
        ChannelMessage t;
        t <- mod_3951.get(0);
        mod_3955.put(0, t);
    endrule
    rule rule_5141;
        ChannelMessage t;
        t <- mod_3970.get(1);
        mod_3945.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3937.put(0, t);
        end
        if (i == 1) begin
            mod_3953.put(0, t);
        end
        if (i == 2) begin
            mod_3959.put(0, t);
        end
        if (i == 3) begin
            mod_3967.put(0, t);
        end
        if (i == 4) begin
            mod_3973.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_3941.get(0);
        end
        if (i == 2) begin
            t <- mod_3941.get(1);
        end
        if (i == 1) begin
            t <- mod_3941.get(2);
        end
        if (i == 3) begin
            t <- mod_3953.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6131 (Operation_IFC);
    Operation_IFC mod_3978_inner <- mkReshape(2, 64);
    Operation_IFC mod_3978 <- mkDebugOperation(mod_3978_inner, "mod_3978");
    Operation_IFC mod_3979_inner <- mkFlatten(1);
    Operation_IFC mod_3979 <- mkDebugOperation(mod_3979_inner, "mod_3979");
    Operation_IFC mod_3980_inner <- mkFlatten(2);
    Operation_IFC mod_3980 <- mkDebugOperation(mod_3980_inner, "mod_3980");
    Operation_IFC mod_3981_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_3981 <- mkDebugOperation(mod_3981_inner, "mod_3981");
    Broadcast_IFC#(4) mod_3982_inner <- mkBroadcast(4);
    Operation_IFC mod_3982 <- mkDebugOperation(mod_3982_inner.op, "mod_3982");
    PMU_IFC mod_3983_bufferize <- mkPMU(2);
    Operation_IFC mod_3983_inner = mod_3983_bufferize.operation;
    Operation_IFC mod_3983 <- mkDebugOperation(mod_3983_inner, "mod_3983");
    Broadcast_IFC#(2) mod_3984_inner <- mkBroadcast(2);
    Operation_IFC mod_3984 <- mkDebugOperation(mod_3984_inner.op, "mod_3984");
    PMU_IFC mod_3985_bufferize <- mkPMU(1);
    Operation_IFC mod_3985_inner = mod_3985_bufferize.operation;
    Operation_IFC mod_3985 <- mkDebugOperation(mod_3985_inner, "mod_3985");
    Operation_IFC mod_3986_inner <- mkBinaryMap(1059, matmul_t_tile);
    Operation_IFC mod_3986 <- mkDebugOperation(mod_3986_inner, "mod_3986");
    Operation_IFC mod_3987_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3987 <- mkDebugOperation(mod_3987_inner, "mod_3987");
    Operation_IFC mod_3988_inner <- mkBinaryMap(1827, mul_tile);
    Operation_IFC mod_3988 <- mkDebugOperation(mod_3988_inner, "mod_3988");
    PMU_IFC mod_3989_bufferize <- mkPMU(1);
    Operation_IFC mod_3989_inner = mod_3989_bufferize.operation;
    Operation_IFC mod_3989 <- mkDebugOperation(mod_3989_inner, "mod_3989");
    Operation_IFC mod_3990_inner <- mkBinaryMap(2369, matmul_t_tile);
    Operation_IFC mod_3990 <- mkDebugOperation(mod_3990_inner, "mod_3990");
    Operation_IFC mod_3991_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_3991 <- mkDebugOperation(mod_3991_inner, "mod_3991");
    Operation_IFC mod_3992_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_3992 <- mkDebugOperation(mod_3992_inner, "mod_3992");
    Operation_IFC mod_3993_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_3993 <- mkDebugOperation(mod_3993_inner, "mod_3993");
    Operation_IFC mod_3994_inner <- mkBinaryMap(2726, mul_tile);
    Operation_IFC mod_3994 <- mkDebugOperation(mod_3994_inner, "mod_3994");
    PMU_IFC mod_3995_bufferize <- mkPMU(1);
    Operation_IFC mod_3995_inner = mod_3995_bufferize.operation;
    Operation_IFC mod_3995 <- mkDebugOperation(mod_3995_inner, "mod_3995");
    PMU_IFC mod_3996_bufferize <- mkPMU(2);
    Operation_IFC mod_3996_inner = mod_3996_bufferize.operation;
    Operation_IFC mod_3996 <- mkDebugOperation(mod_3996_inner, "mod_3996");
    PMU_IFC mod_3997_bufferize <- mkPMU(2);
    Operation_IFC mod_3997_inner = mod_3997_bufferize.operation;
    Operation_IFC mod_3997 <- mkDebugOperation(mod_3997_inner, "mod_3997");
    Operation_IFC mod_3998_inner <- mkRepeatStatic(8);
    Operation_IFC mod_3998 <- mkDebugOperation(mod_3998_inner, "mod_3998");
    Operation_IFC mod_3999_inner <- mkFlatten(1);
    Operation_IFC mod_3999 <- mkDebugOperation(mod_3999_inner, "mod_3999");
    Operation_IFC mod_4000_inner <- mkFlatten(0);
    Operation_IFC mod_4000 <- mkDebugOperation(mod_4000_inner, "mod_4000");
    Operation_IFC mod_4001_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4001 <- mkDebugOperation(mod_4001_inner, "mod_4001");
    Operation_IFC mod_4002_inner <- mkUnaryMap(1699, silu_tile);
    Operation_IFC mod_4002 <- mkDebugOperation(mod_4002_inner, "mod_4002");
    Operation_IFC mod_4003_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4003 <- mkDebugOperation(mod_4003_inner, "mod_4003");
    Operation_IFC mod_4004_inner <- mkBinaryMap(1571, matmul_t_tile);
    Operation_IFC mod_4004 <- mkDebugOperation(mod_4004_inner, "mod_4004");
    PMU_IFC mod_4005_bufferize <- mkPMU(2);
    Operation_IFC mod_4005_inner = mod_4005_bufferize.operation;
    Operation_IFC mod_4005 <- mkDebugOperation(mod_4005_inner, "mod_4005");
    Operation_IFC mod_4006_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4006 <- mkDebugOperation(mod_4006_inner, "mod_4006");
    Operation_IFC mod_4007_inner <- mkFlatten(1);
    Operation_IFC mod_4007 <- mkDebugOperation(mod_4007_inner, "mod_4007");
    Operation_IFC mod_4008_inner <- mkFlatten(0);
    Operation_IFC mod_4008 <- mkDebugOperation(mod_4008_inner, "mod_4008");
    PMU_IFC mod_4009_bufferize <- mkPMU(1);
    Operation_IFC mod_4009_inner = mod_4009_bufferize.operation;
    Operation_IFC mod_4009 <- mkDebugOperation(mod_4009_inner, "mod_4009");
    Operation_IFC mod_4010_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4010 <- mkDebugOperation(mod_4010_inner, "mod_4010");
    PMU_IFC mod_4011_bufferize <- mkPMU(2);
    Operation_IFC mod_4011_inner = mod_4011_bufferize.operation;
    Operation_IFC mod_4011 <- mkDebugOperation(mod_4011_inner, "mod_4011");
    Operation_IFC mod_4012_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4012 <- mkDebugOperation(mod_4012_inner, "mod_4012");
    Operation_IFC mod_4013_inner <- mkFlatten(1);
    Operation_IFC mod_4013 <- mkDebugOperation(mod_4013_inner, "mod_4013");
    Operation_IFC mod_4014_inner <- mkFlatten(0);
    Operation_IFC mod_4014 <- mkDebugOperation(mod_4014_inner, "mod_4014");
    Operation_IFC mod_4015_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4015 <- mkDebugOperation(mod_4015_inner, "mod_4015");
    Operation_IFC mod_4016_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4016 <- mkDebugOperation(mod_4016_inner, "mod_4016");
    PMU_IFC mod_4017_bufferize <- mkPMU(2);
    Operation_IFC mod_4017_inner = mod_4017_bufferize.operation;
    Operation_IFC mod_4017 <- mkDebugOperation(mod_4017_inner, "mod_4017");
    rule rule_5142;
        ChannelMessage t;
        t <- mod_3985.get(1);
        mod_3986.put(0, t);
    endrule
    rule rule_5143;
        ChannelMessage t;
        t <- mod_4017.get(0);
        mod_4017.put(1, t);
    endrule
    rule rule_5144;
        ChannelMessage t;
        t <- mod_3997.get(0);
        mod_3998.put(0, t);
    endrule
    rule rule_5145;
        ChannelMessage t;
        t <- mod_3993.get(1);
        mod_3994.put(1, t);
    endrule
    rule rule_5146;
        ChannelMessage t;
        t <- mod_4011.get(1);
        mod_3986.put(1, t);
    endrule
    rule rule_5147;
        ChannelMessage t;
        t <- mod_3981.get(1);
        mod_3982.put(0, t);
    endrule
    rule rule_5148;
        ChannelMessage t;
        t <- mod_4010.get(0);
        mod_4009.put(1, t);
    endrule
    rule rule_5149;
        ChannelMessage t;
        t <- mod_3984.get(1);
        mod_3985.put(0, t);
    endrule
    rule rule_5150;
        ChannelMessage t;
        t <- mod_3980.get(0);
        mod_3981.put(0, t);
    endrule
    rule rule_5151;
        ChannelMessage t;
        t <- mod_4008.get(0);
        mod_4007.put(0, t);
    endrule
    rule rule_5152;
        ChannelMessage t;
        t <- mod_4007.get(0);
        mod_4005.put(0, t);
    endrule
    rule rule_5153;
        ChannelMessage t;
        t <- mod_3996.get(0);
        mod_3996.put(1, t);
    endrule
    rule rule_5154;
        ChannelMessage t;
        t <- mod_4017.get(1);
        mod_3981.put(1, t);
    endrule
    rule rule_5155;
        ChannelMessage t;
        t <- mod_3995.get(0);
        mod_3995.put(1, t);
    endrule
    rule rule_5156;
        ChannelMessage t;
        t <- mod_3987.get(0);
        mod_3988.put(0, t);
    endrule
    rule rule_5157;
        ChannelMessage t;
        t <- mod_3988.get(0);
        mod_3989.put(0, t);
    endrule
    rule rule_5158;
        ChannelMessage t;
        t <- mod_3993.get(0);
        mod_3995.put(0, t);
    endrule
    rule rule_5159;
        ChannelMessage t;
        t <- mod_3995.get(1);
        mod_3993.put(1, t);
    endrule
    rule rule_5160;
        ChannelMessage t;
        t <- mod_3999.get(0);
        mod_3997.put(0, t);
    endrule
    rule rule_5161;
        ChannelMessage t;
        t <- mod_3989.get(0);
        mod_4001.put(0, t);
    endrule
    rule rule_5162;
        ChannelMessage t;
        t <- mod_4014.get(0);
        mod_4013.put(0, t);
    endrule
    rule rule_5163;
        ChannelMessage t;
        t <- mod_3978.get(0);
        mod_3979.put(0, t);
    endrule
    rule rule_5164;
        ChannelMessage t;
        t <- mod_3982.get(3);
        mod_3983.put(0, t);
    endrule
    rule rule_5165;
        ChannelMessage t;
        t <- mod_3991.get(0);
        mod_3992.put(0, t);
    endrule
    rule rule_5166;
        ChannelMessage t;
        t <- mod_4005.get(0);
        mod_4006.put(0, t);
    endrule
    rule rule_5167;
        ChannelMessage t;
        t <- mod_4006.get(0);
        mod_4005.put(1, t);
    endrule
    rule rule_5168;
        ChannelMessage t;
        t <- mod_4000.get(0);
        mod_3999.put(0, t);
    endrule
    rule rule_5169;
        ChannelMessage t;
        t <- mod_4005.get(1);
        mod_4004.put(1, t);
    endrule
    rule rule_5170;
        ChannelMessage t;
        t <- mod_3984.get(0);
        mod_4009.put(0, t);
    endrule
    rule rule_5171;
        ChannelMessage t;
        t <- mod_4013.get(0);
        mod_4011.put(0, t);
    endrule
    rule rule_5172;
        ChannelMessage t;
        t <- mod_3996.get(1);
        mod_3992.put(1, t);
    endrule
    rule rule_5173;
        ChannelMessage t;
        t <- mod_4002.get(0);
        mod_3988.put(1, t);
    endrule
    rule rule_5174;
        ChannelMessage t;
        t <- mod_4009.get(1);
        mod_4004.put(0, t);
    endrule
    rule rule_5175;
        ChannelMessage t;
        t <- mod_3983.get(0);
        mod_4016.put(0, t);
    endrule
    rule rule_5176;
        ChannelMessage t;
        t <- mod_3986.get(0);
        mod_3987.put(0, t);
    endrule
    rule rule_5177;
        ChannelMessage t;
        t <- mod_3985.get(0);
        mod_4015.put(0, t);
    endrule
    rule rule_5178;
        ChannelMessage t;
        t <- mod_4011.get(0);
        mod_4012.put(0, t);
    endrule
    rule rule_5179;
        ChannelMessage t;
        t <- mod_4012.get(0);
        mod_4011.put(1, t);
    endrule
    rule rule_5180;
        ChannelMessage t;
        t <- mod_3997.get(1);
        mod_3990.put(1, t);
    endrule
    rule rule_5181;
        ChannelMessage t;
        t <- mod_4001.get(0);
        mod_3989.put(1, t);
    endrule
    rule rule_5182;
        ChannelMessage t;
        t <- mod_3979.get(0);
        mod_3980.put(0, t);
    endrule
    rule rule_5183;
        ChannelMessage t;
        t <- mod_4003.get(0);
        mod_4002.put(0, t);
    endrule
    rule rule_5184;
        ChannelMessage t;
        t <- mod_4009.get(0);
        mod_4010.put(0, t);
    endrule
    rule rule_5185;
        ChannelMessage t;
        t <- mod_4015.get(0);
        mod_3985.put(1, t);
    endrule
    rule rule_5186;
        ChannelMessage t;
        t <- mod_3990.get(0);
        mod_3991.put(0, t);
    endrule
    rule rule_5187;
        ChannelMessage t;
        t <- mod_3992.get(1);
        mod_3993.put(0, t);
    endrule
    rule rule_5188;
        ChannelMessage t;
        t <- mod_3983.get(1);
        mod_3984.put(0, t);
    endrule
    rule rule_5189;
        ChannelMessage t;
        t <- mod_3989.get(1);
        mod_3990.put(0, t);
    endrule
    rule rule_5190;
        ChannelMessage t;
        t <- mod_4004.get(0);
        mod_4003.put(0, t);
    endrule
    rule rule_5191;
        ChannelMessage t;
        t <- mod_3981.get(0);
        mod_4017.put(0, t);
    endrule
    rule rule_5192;
        ChannelMessage t;
        t <- mod_3998.get(0);
        mod_3997.put(1, t);
    endrule
    rule rule_5193;
        ChannelMessage t;
        t <- mod_4016.get(0);
        mod_3983.put(1, t);
    endrule
    rule rule_5194;
        ChannelMessage t;
        t <- mod_3992.get(0);
        mod_3996.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_3978.put(0, t);
        end
        if (i == 1) begin
            mod_3994.put(0, t);
        end
        if (i == 2) begin
            mod_4000.put(0, t);
        end
        if (i == 3) begin
            mod_4008.put(0, t);
        end
        if (i == 4) begin
            mod_4014.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_3982.get(0);
        end
        if (i == 2) begin
            t <- mod_3982.get(1);
        end
        if (i == 3) begin
            t <- mod_3982.get(2);
        end
        if (i == 0) begin
            t <- mod_3994.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6132 (Operation_IFC);
    Operation_IFC mod_4019_inner <- mkReshape(2, 64);
    Operation_IFC mod_4019 <- mkDebugOperation(mod_4019_inner, "mod_4019");
    Operation_IFC mod_4020_inner <- mkFlatten(1);
    Operation_IFC mod_4020 <- mkDebugOperation(mod_4020_inner, "mod_4020");
    Operation_IFC mod_4021_inner <- mkFlatten(2);
    Operation_IFC mod_4021 <- mkDebugOperation(mod_4021_inner, "mod_4021");
    Operation_IFC mod_4022_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4022 <- mkDebugOperation(mod_4022_inner, "mod_4022");
    Broadcast_IFC#(4) mod_4023_inner <- mkBroadcast(4);
    Operation_IFC mod_4023 <- mkDebugOperation(mod_4023_inner.op, "mod_4023");
    PMU_IFC mod_4024_bufferize <- mkPMU(2);
    Operation_IFC mod_4024_inner = mod_4024_bufferize.operation;
    Operation_IFC mod_4024 <- mkDebugOperation(mod_4024_inner, "mod_4024");
    Broadcast_IFC#(2) mod_4025_inner <- mkBroadcast(2);
    Operation_IFC mod_4025 <- mkDebugOperation(mod_4025_inner.op, "mod_4025");
    PMU_IFC mod_4026_bufferize <- mkPMU(1);
    Operation_IFC mod_4026_inner = mod_4026_bufferize.operation;
    Operation_IFC mod_4026 <- mkDebugOperation(mod_4026_inner, "mod_4026");
    Operation_IFC mod_4027_inner <- mkBinaryMap(1058, matmul_t_tile);
    Operation_IFC mod_4027 <- mkDebugOperation(mod_4027_inner, "mod_4027");
    Operation_IFC mod_4028_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4028 <- mkDebugOperation(mod_4028_inner, "mod_4028");
    Operation_IFC mod_4029_inner <- mkBinaryMap(1826, mul_tile);
    Operation_IFC mod_4029 <- mkDebugOperation(mod_4029_inner, "mod_4029");
    PMU_IFC mod_4030_bufferize <- mkPMU(1);
    Operation_IFC mod_4030_inner = mod_4030_bufferize.operation;
    Operation_IFC mod_4030 <- mkDebugOperation(mod_4030_inner, "mod_4030");
    Operation_IFC mod_4031_inner <- mkBinaryMap(2367, matmul_t_tile);
    Operation_IFC mod_4031 <- mkDebugOperation(mod_4031_inner, "mod_4031");
    Operation_IFC mod_4032_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4032 <- mkDebugOperation(mod_4032_inner, "mod_4032");
    Operation_IFC mod_4033_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4033 <- mkDebugOperation(mod_4033_inner, "mod_4033");
    Operation_IFC mod_4034_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4034 <- mkDebugOperation(mod_4034_inner, "mod_4034");
    Operation_IFC mod_4035_inner <- mkBinaryMap(2725, mul_tile);
    Operation_IFC mod_4035 <- mkDebugOperation(mod_4035_inner, "mod_4035");
    PMU_IFC mod_4036_bufferize <- mkPMU(1);
    Operation_IFC mod_4036_inner = mod_4036_bufferize.operation;
    Operation_IFC mod_4036 <- mkDebugOperation(mod_4036_inner, "mod_4036");
    PMU_IFC mod_4037_bufferize <- mkPMU(2);
    Operation_IFC mod_4037_inner = mod_4037_bufferize.operation;
    Operation_IFC mod_4037 <- mkDebugOperation(mod_4037_inner, "mod_4037");
    PMU_IFC mod_4038_bufferize <- mkPMU(2);
    Operation_IFC mod_4038_inner = mod_4038_bufferize.operation;
    Operation_IFC mod_4038 <- mkDebugOperation(mod_4038_inner, "mod_4038");
    Operation_IFC mod_4039_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4039 <- mkDebugOperation(mod_4039_inner, "mod_4039");
    Operation_IFC mod_4040_inner <- mkFlatten(1);
    Operation_IFC mod_4040 <- mkDebugOperation(mod_4040_inner, "mod_4040");
    Operation_IFC mod_4041_inner <- mkFlatten(0);
    Operation_IFC mod_4041 <- mkDebugOperation(mod_4041_inner, "mod_4041");
    Operation_IFC mod_4042_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4042 <- mkDebugOperation(mod_4042_inner, "mod_4042");
    Operation_IFC mod_4043_inner <- mkUnaryMap(1698, silu_tile);
    Operation_IFC mod_4043 <- mkDebugOperation(mod_4043_inner, "mod_4043");
    Operation_IFC mod_4044_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4044 <- mkDebugOperation(mod_4044_inner, "mod_4044");
    Operation_IFC mod_4045_inner <- mkBinaryMap(1570, matmul_t_tile);
    Operation_IFC mod_4045 <- mkDebugOperation(mod_4045_inner, "mod_4045");
    PMU_IFC mod_4046_bufferize <- mkPMU(2);
    Operation_IFC mod_4046_inner = mod_4046_bufferize.operation;
    Operation_IFC mod_4046 <- mkDebugOperation(mod_4046_inner, "mod_4046");
    Operation_IFC mod_4047_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4047 <- mkDebugOperation(mod_4047_inner, "mod_4047");
    Operation_IFC mod_4048_inner <- mkFlatten(1);
    Operation_IFC mod_4048 <- mkDebugOperation(mod_4048_inner, "mod_4048");
    Operation_IFC mod_4049_inner <- mkFlatten(0);
    Operation_IFC mod_4049 <- mkDebugOperation(mod_4049_inner, "mod_4049");
    PMU_IFC mod_4050_bufferize <- mkPMU(1);
    Operation_IFC mod_4050_inner = mod_4050_bufferize.operation;
    Operation_IFC mod_4050 <- mkDebugOperation(mod_4050_inner, "mod_4050");
    Operation_IFC mod_4051_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4051 <- mkDebugOperation(mod_4051_inner, "mod_4051");
    PMU_IFC mod_4052_bufferize <- mkPMU(2);
    Operation_IFC mod_4052_inner = mod_4052_bufferize.operation;
    Operation_IFC mod_4052 <- mkDebugOperation(mod_4052_inner, "mod_4052");
    Operation_IFC mod_4053_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4053 <- mkDebugOperation(mod_4053_inner, "mod_4053");
    Operation_IFC mod_4054_inner <- mkFlatten(1);
    Operation_IFC mod_4054 <- mkDebugOperation(mod_4054_inner, "mod_4054");
    Operation_IFC mod_4055_inner <- mkFlatten(0);
    Operation_IFC mod_4055 <- mkDebugOperation(mod_4055_inner, "mod_4055");
    Operation_IFC mod_4056_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4056 <- mkDebugOperation(mod_4056_inner, "mod_4056");
    Operation_IFC mod_4057_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4057 <- mkDebugOperation(mod_4057_inner, "mod_4057");
    PMU_IFC mod_4058_bufferize <- mkPMU(2);
    Operation_IFC mod_4058_inner = mod_4058_bufferize.operation;
    Operation_IFC mod_4058 <- mkDebugOperation(mod_4058_inner, "mod_4058");
    rule rule_5195;
        ChannelMessage t;
        t <- mod_4026.get(1);
        mod_4027.put(0, t);
    endrule
    rule rule_5196;
        ChannelMessage t;
        t <- mod_4037.get(0);
        mod_4037.put(1, t);
    endrule
    rule rule_5197;
        ChannelMessage t;
        t <- mod_4019.get(0);
        mod_4020.put(0, t);
    endrule
    rule rule_5198;
        ChannelMessage t;
        t <- mod_4034.get(0);
        mod_4036.put(0, t);
    endrule
    rule rule_5199;
        ChannelMessage t;
        t <- mod_4033.get(1);
        mod_4034.put(0, t);
    endrule
    rule rule_5200;
        ChannelMessage t;
        t <- mod_4036.get(1);
        mod_4034.put(1, t);
    endrule
    rule rule_5201;
        ChannelMessage t;
        t <- mod_4046.get(1);
        mod_4045.put(1, t);
    endrule
    rule rule_5202;
        ChannelMessage t;
        t <- mod_4058.get(1);
        mod_4022.put(1, t);
    endrule
    rule rule_5203;
        ChannelMessage t;
        t <- mod_4042.get(0);
        mod_4030.put(1, t);
    endrule
    rule rule_5204;
        ChannelMessage t;
        t <- mod_4052.get(0);
        mod_4053.put(0, t);
    endrule
    rule rule_5205;
        ChannelMessage t;
        t <- mod_4054.get(0);
        mod_4052.put(0, t);
    endrule
    rule rule_5206;
        ChannelMessage t;
        t <- mod_4023.get(3);
        mod_4024.put(0, t);
    endrule
    rule rule_5207;
        ChannelMessage t;
        t <- mod_4040.get(0);
        mod_4038.put(0, t);
    endrule
    rule rule_5208;
        ChannelMessage t;
        t <- mod_4051.get(0);
        mod_4050.put(1, t);
    endrule
    rule rule_5209;
        ChannelMessage t;
        t <- mod_4038.get(1);
        mod_4031.put(1, t);
    endrule
    rule rule_5210;
        ChannelMessage t;
        t <- mod_4022.get(0);
        mod_4058.put(0, t);
    endrule
    rule rule_5211;
        ChannelMessage t;
        t <- mod_4056.get(0);
        mod_4026.put(1, t);
    endrule
    rule rule_5212;
        ChannelMessage t;
        t <- mod_4050.get(0);
        mod_4051.put(0, t);
    endrule
    rule rule_5213;
        ChannelMessage t;
        t <- mod_4032.get(0);
        mod_4033.put(0, t);
    endrule
    rule rule_5214;
        ChannelMessage t;
        t <- mod_4031.get(0);
        mod_4032.put(0, t);
    endrule
    rule rule_5215;
        ChannelMessage t;
        t <- mod_4034.get(1);
        mod_4035.put(1, t);
    endrule
    rule rule_5216;
        ChannelMessage t;
        t <- mod_4022.get(1);
        mod_4023.put(0, t);
    endrule
    rule rule_5217;
        ChannelMessage t;
        t <- mod_4030.get(0);
        mod_4042.put(0, t);
    endrule
    rule rule_5218;
        ChannelMessage t;
        t <- mod_4043.get(0);
        mod_4029.put(1, t);
    endrule
    rule rule_5219;
        ChannelMessage t;
        t <- mod_4039.get(0);
        mod_4038.put(1, t);
    endrule
    rule rule_5220;
        ChannelMessage t;
        t <- mod_4028.get(0);
        mod_4029.put(0, t);
    endrule
    rule rule_5221;
        ChannelMessage t;
        t <- mod_4045.get(0);
        mod_4044.put(0, t);
    endrule
    rule rule_5222;
        ChannelMessage t;
        t <- mod_4052.get(1);
        mod_4027.put(1, t);
    endrule
    rule rule_5223;
        ChannelMessage t;
        t <- mod_4038.get(0);
        mod_4039.put(0, t);
    endrule
    rule rule_5224;
        ChannelMessage t;
        t <- mod_4024.get(1);
        mod_4025.put(0, t);
    endrule
    rule rule_5225;
        ChannelMessage t;
        t <- mod_4026.get(0);
        mod_4056.put(0, t);
    endrule
    rule rule_5226;
        ChannelMessage t;
        t <- mod_4020.get(0);
        mod_4021.put(0, t);
    endrule
    rule rule_5227;
        ChannelMessage t;
        t <- mod_4033.get(0);
        mod_4037.put(0, t);
    endrule
    rule rule_5228;
        ChannelMessage t;
        t <- mod_4036.get(0);
        mod_4036.put(1, t);
    endrule
    rule rule_5229;
        ChannelMessage t;
        t <- mod_4030.get(1);
        mod_4031.put(0, t);
    endrule
    rule rule_5230;
        ChannelMessage t;
        t <- mod_4041.get(0);
        mod_4040.put(0, t);
    endrule
    rule rule_5231;
        ChannelMessage t;
        t <- mod_4027.get(0);
        mod_4028.put(0, t);
    endrule
    rule rule_5232;
        ChannelMessage t;
        t <- mod_4058.get(0);
        mod_4058.put(1, t);
    endrule
    rule rule_5233;
        ChannelMessage t;
        t <- mod_4025.get(1);
        mod_4026.put(0, t);
    endrule
    rule rule_5234;
        ChannelMessage t;
        t <- mod_4048.get(0);
        mod_4046.put(0, t);
    endrule
    rule rule_5235;
        ChannelMessage t;
        t <- mod_4047.get(0);
        mod_4046.put(1, t);
    endrule
    rule rule_5236;
        ChannelMessage t;
        t <- mod_4055.get(0);
        mod_4054.put(0, t);
    endrule
    rule rule_5237;
        ChannelMessage t;
        t <- mod_4025.get(0);
        mod_4050.put(0, t);
    endrule
    rule rule_5238;
        ChannelMessage t;
        t <- mod_4044.get(0);
        mod_4043.put(0, t);
    endrule
    rule rule_5239;
        ChannelMessage t;
        t <- mod_4029.get(0);
        mod_4030.put(0, t);
    endrule
    rule rule_5240;
        ChannelMessage t;
        t <- mod_4053.get(0);
        mod_4052.put(1, t);
    endrule
    rule rule_5241;
        ChannelMessage t;
        t <- mod_4037.get(1);
        mod_4033.put(1, t);
    endrule
    rule rule_5242;
        ChannelMessage t;
        t <- mod_4049.get(0);
        mod_4048.put(0, t);
    endrule
    rule rule_5243;
        ChannelMessage t;
        t <- mod_4024.get(0);
        mod_4057.put(0, t);
    endrule
    rule rule_5244;
        ChannelMessage t;
        t <- mod_4050.get(1);
        mod_4045.put(0, t);
    endrule
    rule rule_5245;
        ChannelMessage t;
        t <- mod_4057.get(0);
        mod_4024.put(1, t);
    endrule
    rule rule_5246;
        ChannelMessage t;
        t <- mod_4021.get(0);
        mod_4022.put(0, t);
    endrule
    rule rule_5247;
        ChannelMessage t;
        t <- mod_4046.get(0);
        mod_4047.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4019.put(0, t);
        end
        if (i == 1) begin
            mod_4035.put(0, t);
        end
        if (i == 2) begin
            mod_4041.put(0, t);
        end
        if (i == 3) begin
            mod_4049.put(0, t);
        end
        if (i == 4) begin
            mod_4055.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_4023.get(0);
        end
        if (i == 2) begin
            t <- mod_4023.get(1);
        end
        if (i == 0) begin
            t <- mod_4023.get(2);
        end
        if (i == 1) begin
            t <- mod_4035.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6133 (Operation_IFC);
    Operation_IFC mod_4060_inner <- mkReshape(2, 64);
    Operation_IFC mod_4060 <- mkDebugOperation(mod_4060_inner, "mod_4060");
    Operation_IFC mod_4061_inner <- mkFlatten(1);
    Operation_IFC mod_4061 <- mkDebugOperation(mod_4061_inner, "mod_4061");
    Operation_IFC mod_4062_inner <- mkFlatten(2);
    Operation_IFC mod_4062 <- mkDebugOperation(mod_4062_inner, "mod_4062");
    Operation_IFC mod_4063_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4063 <- mkDebugOperation(mod_4063_inner, "mod_4063");
    Broadcast_IFC#(4) mod_4064_inner <- mkBroadcast(4);
    Operation_IFC mod_4064 <- mkDebugOperation(mod_4064_inner.op, "mod_4064");
    PMU_IFC mod_4065_bufferize <- mkPMU(2);
    Operation_IFC mod_4065_inner = mod_4065_bufferize.operation;
    Operation_IFC mod_4065 <- mkDebugOperation(mod_4065_inner, "mod_4065");
    Broadcast_IFC#(2) mod_4066_inner <- mkBroadcast(2);
    Operation_IFC mod_4066 <- mkDebugOperation(mod_4066_inner.op, "mod_4066");
    PMU_IFC mod_4067_bufferize <- mkPMU(1);
    Operation_IFC mod_4067_inner = mod_4067_bufferize.operation;
    Operation_IFC mod_4067 <- mkDebugOperation(mod_4067_inner, "mod_4067");
    Operation_IFC mod_4068_inner <- mkBinaryMap(1057, matmul_t_tile);
    Operation_IFC mod_4068 <- mkDebugOperation(mod_4068_inner, "mod_4068");
    Operation_IFC mod_4069_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4069 <- mkDebugOperation(mod_4069_inner, "mod_4069");
    Operation_IFC mod_4070_inner <- mkBinaryMap(1825, mul_tile);
    Operation_IFC mod_4070 <- mkDebugOperation(mod_4070_inner, "mod_4070");
    PMU_IFC mod_4071_bufferize <- mkPMU(1);
    Operation_IFC mod_4071_inner = mod_4071_bufferize.operation;
    Operation_IFC mod_4071 <- mkDebugOperation(mod_4071_inner, "mod_4071");
    Operation_IFC mod_4072_inner <- mkBinaryMap(2365, matmul_t_tile);
    Operation_IFC mod_4072 <- mkDebugOperation(mod_4072_inner, "mod_4072");
    Operation_IFC mod_4073_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4073 <- mkDebugOperation(mod_4073_inner, "mod_4073");
    Operation_IFC mod_4074_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4074 <- mkDebugOperation(mod_4074_inner, "mod_4074");
    Operation_IFC mod_4075_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4075 <- mkDebugOperation(mod_4075_inner, "mod_4075");
    Operation_IFC mod_4076_inner <- mkBinaryMap(2724, mul_tile);
    Operation_IFC mod_4076 <- mkDebugOperation(mod_4076_inner, "mod_4076");
    PMU_IFC mod_4077_bufferize <- mkPMU(1);
    Operation_IFC mod_4077_inner = mod_4077_bufferize.operation;
    Operation_IFC mod_4077 <- mkDebugOperation(mod_4077_inner, "mod_4077");
    PMU_IFC mod_4078_bufferize <- mkPMU(2);
    Operation_IFC mod_4078_inner = mod_4078_bufferize.operation;
    Operation_IFC mod_4078 <- mkDebugOperation(mod_4078_inner, "mod_4078");
    PMU_IFC mod_4079_bufferize <- mkPMU(2);
    Operation_IFC mod_4079_inner = mod_4079_bufferize.operation;
    Operation_IFC mod_4079 <- mkDebugOperation(mod_4079_inner, "mod_4079");
    Operation_IFC mod_4080_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4080 <- mkDebugOperation(mod_4080_inner, "mod_4080");
    Operation_IFC mod_4081_inner <- mkFlatten(1);
    Operation_IFC mod_4081 <- mkDebugOperation(mod_4081_inner, "mod_4081");
    Operation_IFC mod_4082_inner <- mkFlatten(0);
    Operation_IFC mod_4082 <- mkDebugOperation(mod_4082_inner, "mod_4082");
    Operation_IFC mod_4083_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4083 <- mkDebugOperation(mod_4083_inner, "mod_4083");
    Operation_IFC mod_4084_inner <- mkUnaryMap(1697, silu_tile);
    Operation_IFC mod_4084 <- mkDebugOperation(mod_4084_inner, "mod_4084");
    Operation_IFC mod_4085_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4085 <- mkDebugOperation(mod_4085_inner, "mod_4085");
    Operation_IFC mod_4086_inner <- mkBinaryMap(1569, matmul_t_tile);
    Operation_IFC mod_4086 <- mkDebugOperation(mod_4086_inner, "mod_4086");
    PMU_IFC mod_4087_bufferize <- mkPMU(2);
    Operation_IFC mod_4087_inner = mod_4087_bufferize.operation;
    Operation_IFC mod_4087 <- mkDebugOperation(mod_4087_inner, "mod_4087");
    Operation_IFC mod_4088_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4088 <- mkDebugOperation(mod_4088_inner, "mod_4088");
    Operation_IFC mod_4089_inner <- mkFlatten(1);
    Operation_IFC mod_4089 <- mkDebugOperation(mod_4089_inner, "mod_4089");
    Operation_IFC mod_4090_inner <- mkFlatten(0);
    Operation_IFC mod_4090 <- mkDebugOperation(mod_4090_inner, "mod_4090");
    PMU_IFC mod_4091_bufferize <- mkPMU(1);
    Operation_IFC mod_4091_inner = mod_4091_bufferize.operation;
    Operation_IFC mod_4091 <- mkDebugOperation(mod_4091_inner, "mod_4091");
    Operation_IFC mod_4092_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4092 <- mkDebugOperation(mod_4092_inner, "mod_4092");
    PMU_IFC mod_4093_bufferize <- mkPMU(2);
    Operation_IFC mod_4093_inner = mod_4093_bufferize.operation;
    Operation_IFC mod_4093 <- mkDebugOperation(mod_4093_inner, "mod_4093");
    Operation_IFC mod_4094_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4094 <- mkDebugOperation(mod_4094_inner, "mod_4094");
    Operation_IFC mod_4095_inner <- mkFlatten(1);
    Operation_IFC mod_4095 <- mkDebugOperation(mod_4095_inner, "mod_4095");
    Operation_IFC mod_4096_inner <- mkFlatten(0);
    Operation_IFC mod_4096 <- mkDebugOperation(mod_4096_inner, "mod_4096");
    Operation_IFC mod_4097_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4097 <- mkDebugOperation(mod_4097_inner, "mod_4097");
    Operation_IFC mod_4098_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4098 <- mkDebugOperation(mod_4098_inner, "mod_4098");
    PMU_IFC mod_4099_bufferize <- mkPMU(2);
    Operation_IFC mod_4099_inner = mod_4099_bufferize.operation;
    Operation_IFC mod_4099 <- mkDebugOperation(mod_4099_inner, "mod_4099");
    rule rule_5248;
        ChannelMessage t;
        t <- mod_4060.get(0);
        mod_4061.put(0, t);
    endrule
    rule rule_5249;
        ChannelMessage t;
        t <- mod_4077.get(0);
        mod_4077.put(1, t);
    endrule
    rule rule_5250;
        ChannelMessage t;
        t <- mod_4064.get(3);
        mod_4065.put(0, t);
    endrule
    rule rule_5251;
        ChannelMessage t;
        t <- mod_4086.get(0);
        mod_4085.put(0, t);
    endrule
    rule rule_5252;
        ChannelMessage t;
        t <- mod_4084.get(0);
        mod_4070.put(1, t);
    endrule
    rule rule_5253;
        ChannelMessage t;
        t <- mod_4073.get(0);
        mod_4074.put(0, t);
    endrule
    rule rule_5254;
        ChannelMessage t;
        t <- mod_4071.get(1);
        mod_4072.put(0, t);
    endrule
    rule rule_5255;
        ChannelMessage t;
        t <- mod_4075.get(0);
        mod_4077.put(0, t);
    endrule
    rule rule_5256;
        ChannelMessage t;
        t <- mod_4070.get(0);
        mod_4071.put(0, t);
    endrule
    rule rule_5257;
        ChannelMessage t;
        t <- mod_4082.get(0);
        mod_4081.put(0, t);
    endrule
    rule rule_5258;
        ChannelMessage t;
        t <- mod_4094.get(0);
        mod_4093.put(1, t);
    endrule
    rule rule_5259;
        ChannelMessage t;
        t <- mod_4092.get(0);
        mod_4091.put(1, t);
    endrule
    rule rule_5260;
        ChannelMessage t;
        t <- mod_4096.get(0);
        mod_4095.put(0, t);
    endrule
    rule rule_5261;
        ChannelMessage t;
        t <- mod_4063.get(0);
        mod_4099.put(0, t);
    endrule
    rule rule_5262;
        ChannelMessage t;
        t <- mod_4098.get(0);
        mod_4065.put(1, t);
    endrule
    rule rule_5263;
        ChannelMessage t;
        t <- mod_4075.get(1);
        mod_4076.put(1, t);
    endrule
    rule rule_5264;
        ChannelMessage t;
        t <- mod_4093.get(1);
        mod_4068.put(1, t);
    endrule
    rule rule_5265;
        ChannelMessage t;
        t <- mod_4091.get(0);
        mod_4092.put(0, t);
    endrule
    rule rule_5266;
        ChannelMessage t;
        t <- mod_4099.get(1);
        mod_4063.put(1, t);
    endrule
    rule rule_5267;
        ChannelMessage t;
        t <- mod_4066.get(0);
        mod_4091.put(0, t);
    endrule
    rule rule_5268;
        ChannelMessage t;
        t <- mod_4085.get(0);
        mod_4084.put(0, t);
    endrule
    rule rule_5269;
        ChannelMessage t;
        t <- mod_4079.get(1);
        mod_4072.put(1, t);
    endrule
    rule rule_5270;
        ChannelMessage t;
        t <- mod_4078.get(0);
        mod_4078.put(1, t);
    endrule
    rule rule_5271;
        ChannelMessage t;
        t <- mod_4080.get(0);
        mod_4079.put(1, t);
    endrule
    rule rule_5272;
        ChannelMessage t;
        t <- mod_4063.get(1);
        mod_4064.put(0, t);
    endrule
    rule rule_5273;
        ChannelMessage t;
        t <- mod_4078.get(1);
        mod_4074.put(1, t);
    endrule
    rule rule_5274;
        ChannelMessage t;
        t <- mod_4071.get(0);
        mod_4083.put(0, t);
    endrule
    rule rule_5275;
        ChannelMessage t;
        t <- mod_4088.get(0);
        mod_4087.put(1, t);
    endrule
    rule rule_5276;
        ChannelMessage t;
        t <- mod_4091.get(1);
        mod_4086.put(0, t);
    endrule
    rule rule_5277;
        ChannelMessage t;
        t <- mod_4097.get(0);
        mod_4067.put(1, t);
    endrule
    rule rule_5278;
        ChannelMessage t;
        t <- mod_4067.get(0);
        mod_4097.put(0, t);
    endrule
    rule rule_5279;
        ChannelMessage t;
        t <- mod_4069.get(0);
        mod_4070.put(0, t);
    endrule
    rule rule_5280;
        ChannelMessage t;
        t <- mod_4066.get(1);
        mod_4067.put(0, t);
    endrule
    rule rule_5281;
        ChannelMessage t;
        t <- mod_4079.get(0);
        mod_4080.put(0, t);
    endrule
    rule rule_5282;
        ChannelMessage t;
        t <- mod_4072.get(0);
        mod_4073.put(0, t);
    endrule
    rule rule_5283;
        ChannelMessage t;
        t <- mod_4087.get(1);
        mod_4086.put(1, t);
    endrule
    rule rule_5284;
        ChannelMessage t;
        t <- mod_4065.get(0);
        mod_4098.put(0, t);
    endrule
    rule rule_5285;
        ChannelMessage t;
        t <- mod_4077.get(1);
        mod_4075.put(1, t);
    endrule
    rule rule_5286;
        ChannelMessage t;
        t <- mod_4068.get(0);
        mod_4069.put(0, t);
    endrule
    rule rule_5287;
        ChannelMessage t;
        t <- mod_4083.get(0);
        mod_4071.put(1, t);
    endrule
    rule rule_5288;
        ChannelMessage t;
        t <- mod_4067.get(1);
        mod_4068.put(0, t);
    endrule
    rule rule_5289;
        ChannelMessage t;
        t <- mod_4089.get(0);
        mod_4087.put(0, t);
    endrule
    rule rule_5290;
        ChannelMessage t;
        t <- mod_4081.get(0);
        mod_4079.put(0, t);
    endrule
    rule rule_5291;
        ChannelMessage t;
        t <- mod_4093.get(0);
        mod_4094.put(0, t);
    endrule
    rule rule_5292;
        ChannelMessage t;
        t <- mod_4074.get(0);
        mod_4078.put(0, t);
    endrule
    rule rule_5293;
        ChannelMessage t;
        t <- mod_4090.get(0);
        mod_4089.put(0, t);
    endrule
    rule rule_5294;
        ChannelMessage t;
        t <- mod_4062.get(0);
        mod_4063.put(0, t);
    endrule
    rule rule_5295;
        ChannelMessage t;
        t <- mod_4074.get(1);
        mod_4075.put(0, t);
    endrule
    rule rule_5296;
        ChannelMessage t;
        t <- mod_4065.get(1);
        mod_4066.put(0, t);
    endrule
    rule rule_5297;
        ChannelMessage t;
        t <- mod_4099.get(0);
        mod_4099.put(1, t);
    endrule
    rule rule_5298;
        ChannelMessage t;
        t <- mod_4095.get(0);
        mod_4093.put(0, t);
    endrule
    rule rule_5299;
        ChannelMessage t;
        t <- mod_4087.get(0);
        mod_4088.put(0, t);
    endrule
    rule rule_5300;
        ChannelMessage t;
        t <- mod_4061.get(0);
        mod_4062.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4060.put(0, t);
        end
        if (i == 1) begin
            mod_4076.put(0, t);
        end
        if (i == 2) begin
            mod_4082.put(0, t);
        end
        if (i == 3) begin
            mod_4090.put(0, t);
        end
        if (i == 4) begin
            mod_4096.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_4064.get(0);
        end
        if (i == 2) begin
            t <- mod_4064.get(1);
        end
        if (i == 0) begin
            t <- mod_4064.get(2);
        end
        if (i == 3) begin
            t <- mod_4076.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6134 (Operation_IFC);
    Operation_IFC mod_4101_inner <- mkReshape(2, 64);
    Operation_IFC mod_4101 <- mkDebugOperation(mod_4101_inner, "mod_4101");
    Operation_IFC mod_4102_inner <- mkFlatten(1);
    Operation_IFC mod_4102 <- mkDebugOperation(mod_4102_inner, "mod_4102");
    Operation_IFC mod_4103_inner <- mkFlatten(2);
    Operation_IFC mod_4103 <- mkDebugOperation(mod_4103_inner, "mod_4103");
    Operation_IFC mod_4104_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4104 <- mkDebugOperation(mod_4104_inner, "mod_4104");
    Broadcast_IFC#(4) mod_4105_inner <- mkBroadcast(4);
    Operation_IFC mod_4105 <- mkDebugOperation(mod_4105_inner.op, "mod_4105");
    PMU_IFC mod_4106_bufferize <- mkPMU(2);
    Operation_IFC mod_4106_inner = mod_4106_bufferize.operation;
    Operation_IFC mod_4106 <- mkDebugOperation(mod_4106_inner, "mod_4106");
    Broadcast_IFC#(2) mod_4107_inner <- mkBroadcast(2);
    Operation_IFC mod_4107 <- mkDebugOperation(mod_4107_inner.op, "mod_4107");
    PMU_IFC mod_4108_bufferize <- mkPMU(1);
    Operation_IFC mod_4108_inner = mod_4108_bufferize.operation;
    Operation_IFC mod_4108 <- mkDebugOperation(mod_4108_inner, "mod_4108");
    Operation_IFC mod_4109_inner <- mkBinaryMap(1056, matmul_t_tile);
    Operation_IFC mod_4109 <- mkDebugOperation(mod_4109_inner, "mod_4109");
    Operation_IFC mod_4110_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4110 <- mkDebugOperation(mod_4110_inner, "mod_4110");
    Operation_IFC mod_4111_inner <- mkBinaryMap(1824, mul_tile);
    Operation_IFC mod_4111 <- mkDebugOperation(mod_4111_inner, "mod_4111");
    PMU_IFC mod_4112_bufferize <- mkPMU(1);
    Operation_IFC mod_4112_inner = mod_4112_bufferize.operation;
    Operation_IFC mod_4112 <- mkDebugOperation(mod_4112_inner, "mod_4112");
    Operation_IFC mod_4113_inner <- mkBinaryMap(2363, matmul_t_tile);
    Operation_IFC mod_4113 <- mkDebugOperation(mod_4113_inner, "mod_4113");
    Operation_IFC mod_4114_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4114 <- mkDebugOperation(mod_4114_inner, "mod_4114");
    Operation_IFC mod_4115_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4115 <- mkDebugOperation(mod_4115_inner, "mod_4115");
    Operation_IFC mod_4116_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4116 <- mkDebugOperation(mod_4116_inner, "mod_4116");
    Operation_IFC mod_4117_inner <- mkBinaryMap(2723, mul_tile);
    Operation_IFC mod_4117 <- mkDebugOperation(mod_4117_inner, "mod_4117");
    PMU_IFC mod_4118_bufferize <- mkPMU(1);
    Operation_IFC mod_4118_inner = mod_4118_bufferize.operation;
    Operation_IFC mod_4118 <- mkDebugOperation(mod_4118_inner, "mod_4118");
    PMU_IFC mod_4119_bufferize <- mkPMU(2);
    Operation_IFC mod_4119_inner = mod_4119_bufferize.operation;
    Operation_IFC mod_4119 <- mkDebugOperation(mod_4119_inner, "mod_4119");
    PMU_IFC mod_4120_bufferize <- mkPMU(2);
    Operation_IFC mod_4120_inner = mod_4120_bufferize.operation;
    Operation_IFC mod_4120 <- mkDebugOperation(mod_4120_inner, "mod_4120");
    Operation_IFC mod_4121_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4121 <- mkDebugOperation(mod_4121_inner, "mod_4121");
    Operation_IFC mod_4122_inner <- mkFlatten(1);
    Operation_IFC mod_4122 <- mkDebugOperation(mod_4122_inner, "mod_4122");
    Operation_IFC mod_4123_inner <- mkFlatten(0);
    Operation_IFC mod_4123 <- mkDebugOperation(mod_4123_inner, "mod_4123");
    Operation_IFC mod_4124_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4124 <- mkDebugOperation(mod_4124_inner, "mod_4124");
    Operation_IFC mod_4125_inner <- mkUnaryMap(1696, silu_tile);
    Operation_IFC mod_4125 <- mkDebugOperation(mod_4125_inner, "mod_4125");
    Operation_IFC mod_4126_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4126 <- mkDebugOperation(mod_4126_inner, "mod_4126");
    Operation_IFC mod_4127_inner <- mkBinaryMap(1568, matmul_t_tile);
    Operation_IFC mod_4127 <- mkDebugOperation(mod_4127_inner, "mod_4127");
    PMU_IFC mod_4128_bufferize <- mkPMU(2);
    Operation_IFC mod_4128_inner = mod_4128_bufferize.operation;
    Operation_IFC mod_4128 <- mkDebugOperation(mod_4128_inner, "mod_4128");
    Operation_IFC mod_4129_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4129 <- mkDebugOperation(mod_4129_inner, "mod_4129");
    Operation_IFC mod_4130_inner <- mkFlatten(1);
    Operation_IFC mod_4130 <- mkDebugOperation(mod_4130_inner, "mod_4130");
    Operation_IFC mod_4131_inner <- mkFlatten(0);
    Operation_IFC mod_4131 <- mkDebugOperation(mod_4131_inner, "mod_4131");
    PMU_IFC mod_4132_bufferize <- mkPMU(1);
    Operation_IFC mod_4132_inner = mod_4132_bufferize.operation;
    Operation_IFC mod_4132 <- mkDebugOperation(mod_4132_inner, "mod_4132");
    Operation_IFC mod_4133_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4133 <- mkDebugOperation(mod_4133_inner, "mod_4133");
    PMU_IFC mod_4134_bufferize <- mkPMU(2);
    Operation_IFC mod_4134_inner = mod_4134_bufferize.operation;
    Operation_IFC mod_4134 <- mkDebugOperation(mod_4134_inner, "mod_4134");
    Operation_IFC mod_4135_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4135 <- mkDebugOperation(mod_4135_inner, "mod_4135");
    Operation_IFC mod_4136_inner <- mkFlatten(1);
    Operation_IFC mod_4136 <- mkDebugOperation(mod_4136_inner, "mod_4136");
    Operation_IFC mod_4137_inner <- mkFlatten(0);
    Operation_IFC mod_4137 <- mkDebugOperation(mod_4137_inner, "mod_4137");
    Operation_IFC mod_4138_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4138 <- mkDebugOperation(mod_4138_inner, "mod_4138");
    Operation_IFC mod_4139_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4139 <- mkDebugOperation(mod_4139_inner, "mod_4139");
    PMU_IFC mod_4140_bufferize <- mkPMU(2);
    Operation_IFC mod_4140_inner = mod_4140_bufferize.operation;
    Operation_IFC mod_4140 <- mkDebugOperation(mod_4140_inner, "mod_4140");
    rule rule_5301;
        ChannelMessage t;
        t <- mod_4137.get(0);
        mod_4136.put(0, t);
    endrule
    rule rule_5302;
        ChannelMessage t;
        t <- mod_4114.get(0);
        mod_4115.put(0, t);
    endrule
    rule rule_5303;
        ChannelMessage t;
        t <- mod_4108.get(0);
        mod_4138.put(0, t);
    endrule
    rule rule_5304;
        ChannelMessage t;
        t <- mod_4133.get(0);
        mod_4132.put(1, t);
    endrule
    rule rule_5305;
        ChannelMessage t;
        t <- mod_4131.get(0);
        mod_4130.put(0, t);
    endrule
    rule rule_5306;
        ChannelMessage t;
        t <- mod_4119.get(1);
        mod_4115.put(1, t);
    endrule
    rule rule_5307;
        ChannelMessage t;
        t <- mod_4102.get(0);
        mod_4103.put(0, t);
    endrule
    rule rule_5308;
        ChannelMessage t;
        t <- mod_4105.get(3);
        mod_4106.put(0, t);
    endrule
    rule rule_5309;
        ChannelMessage t;
        t <- mod_4132.get(1);
        mod_4127.put(0, t);
    endrule
    rule rule_5310;
        ChannelMessage t;
        t <- mod_4107.get(0);
        mod_4132.put(0, t);
    endrule
    rule rule_5311;
        ChannelMessage t;
        t <- mod_4106.get(1);
        mod_4107.put(0, t);
    endrule
    rule rule_5312;
        ChannelMessage t;
        t <- mod_4130.get(0);
        mod_4128.put(0, t);
    endrule
    rule rule_5313;
        ChannelMessage t;
        t <- mod_4128.get(1);
        mod_4127.put(1, t);
    endrule
    rule rule_5314;
        ChannelMessage t;
        t <- mod_4116.get(1);
        mod_4117.put(1, t);
    endrule
    rule rule_5315;
        ChannelMessage t;
        t <- mod_4120.get(0);
        mod_4121.put(0, t);
    endrule
    rule rule_5316;
        ChannelMessage t;
        t <- mod_4128.get(0);
        mod_4129.put(0, t);
    endrule
    rule rule_5317;
        ChannelMessage t;
        t <- mod_4103.get(0);
        mod_4104.put(0, t);
    endrule
    rule rule_5318;
        ChannelMessage t;
        t <- mod_4113.get(0);
        mod_4114.put(0, t);
    endrule
    rule rule_5319;
        ChannelMessage t;
        t <- mod_4127.get(0);
        mod_4126.put(0, t);
    endrule
    rule rule_5320;
        ChannelMessage t;
        t <- mod_4136.get(0);
        mod_4134.put(0, t);
    endrule
    rule rule_5321;
        ChannelMessage t;
        t <- mod_4110.get(0);
        mod_4111.put(0, t);
    endrule
    rule rule_5322;
        ChannelMessage t;
        t <- mod_4112.get(1);
        mod_4113.put(0, t);
    endrule
    rule rule_5323;
        ChannelMessage t;
        t <- mod_4116.get(0);
        mod_4118.put(0, t);
    endrule
    rule rule_5324;
        ChannelMessage t;
        t <- mod_4118.get(0);
        mod_4118.put(1, t);
    endrule
    rule rule_5325;
        ChannelMessage t;
        t <- mod_4118.get(1);
        mod_4116.put(1, t);
    endrule
    rule rule_5326;
        ChannelMessage t;
        t <- mod_4121.get(0);
        mod_4120.put(1, t);
    endrule
    rule rule_5327;
        ChannelMessage t;
        t <- mod_4123.get(0);
        mod_4122.put(0, t);
    endrule
    rule rule_5328;
        ChannelMessage t;
        t <- mod_4134.get(1);
        mod_4109.put(1, t);
    endrule
    rule rule_5329;
        ChannelMessage t;
        t <- mod_4126.get(0);
        mod_4125.put(0, t);
    endrule
    rule rule_5330;
        ChannelMessage t;
        t <- mod_4134.get(0);
        mod_4135.put(0, t);
    endrule
    rule rule_5331;
        ChannelMessage t;
        t <- mod_4140.get(0);
        mod_4140.put(1, t);
    endrule
    rule rule_5332;
        ChannelMessage t;
        t <- mod_4104.get(0);
        mod_4140.put(0, t);
    endrule
    rule rule_5333;
        ChannelMessage t;
        t <- mod_4122.get(0);
        mod_4120.put(0, t);
    endrule
    rule rule_5334;
        ChannelMessage t;
        t <- mod_4112.get(0);
        mod_4124.put(0, t);
    endrule
    rule rule_5335;
        ChannelMessage t;
        t <- mod_4104.get(1);
        mod_4105.put(0, t);
    endrule
    rule rule_5336;
        ChannelMessage t;
        t <- mod_4138.get(0);
        mod_4108.put(1, t);
    endrule
    rule rule_5337;
        ChannelMessage t;
        t <- mod_4119.get(0);
        mod_4119.put(1, t);
    endrule
    rule rule_5338;
        ChannelMessage t;
        t <- mod_4101.get(0);
        mod_4102.put(0, t);
    endrule
    rule rule_5339;
        ChannelMessage t;
        t <- mod_4120.get(1);
        mod_4113.put(1, t);
    endrule
    rule rule_5340;
        ChannelMessage t;
        t <- mod_4115.get(1);
        mod_4116.put(0, t);
    endrule
    rule rule_5341;
        ChannelMessage t;
        t <- mod_4132.get(0);
        mod_4133.put(0, t);
    endrule
    rule rule_5342;
        ChannelMessage t;
        t <- mod_4108.get(1);
        mod_4109.put(0, t);
    endrule
    rule rule_5343;
        ChannelMessage t;
        t <- mod_4107.get(1);
        mod_4108.put(0, t);
    endrule
    rule rule_5344;
        ChannelMessage t;
        t <- mod_4106.get(0);
        mod_4139.put(0, t);
    endrule
    rule rule_5345;
        ChannelMessage t;
        t <- mod_4109.get(0);
        mod_4110.put(0, t);
    endrule
    rule rule_5346;
        ChannelMessage t;
        t <- mod_4115.get(0);
        mod_4119.put(0, t);
    endrule
    rule rule_5347;
        ChannelMessage t;
        t <- mod_4111.get(0);
        mod_4112.put(0, t);
    endrule
    rule rule_5348;
        ChannelMessage t;
        t <- mod_4125.get(0);
        mod_4111.put(1, t);
    endrule
    rule rule_5349;
        ChannelMessage t;
        t <- mod_4129.get(0);
        mod_4128.put(1, t);
    endrule
    rule rule_5350;
        ChannelMessage t;
        t <- mod_4139.get(0);
        mod_4106.put(1, t);
    endrule
    rule rule_5351;
        ChannelMessage t;
        t <- mod_4135.get(0);
        mod_4134.put(1, t);
    endrule
    rule rule_5352;
        ChannelMessage t;
        t <- mod_4140.get(1);
        mod_4104.put(1, t);
    endrule
    rule rule_5353;
        ChannelMessage t;
        t <- mod_4124.get(0);
        mod_4112.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4101.put(0, t);
        end
        if (i == 1) begin
            mod_4117.put(0, t);
        end
        if (i == 2) begin
            mod_4123.put(0, t);
        end
        if (i == 3) begin
            mod_4131.put(0, t);
        end
        if (i == 4) begin
            mod_4137.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_4105.get(0);
        end
        if (i == 0) begin
            t <- mod_4105.get(1);
        end
        if (i == 1) begin
            t <- mod_4105.get(2);
        end
        if (i == 2) begin
            t <- mod_4117.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6135 (Operation_IFC);
    Operation_IFC mod_4142_inner <- mkReshape(2, 64);
    Operation_IFC mod_4142 <- mkDebugOperation(mod_4142_inner, "mod_4142");
    Operation_IFC mod_4143_inner <- mkFlatten(1);
    Operation_IFC mod_4143 <- mkDebugOperation(mod_4143_inner, "mod_4143");
    Operation_IFC mod_4144_inner <- mkFlatten(2);
    Operation_IFC mod_4144 <- mkDebugOperation(mod_4144_inner, "mod_4144");
    Operation_IFC mod_4145_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4145 <- mkDebugOperation(mod_4145_inner, "mod_4145");
    Broadcast_IFC#(4) mod_4146_inner <- mkBroadcast(4);
    Operation_IFC mod_4146 <- mkDebugOperation(mod_4146_inner.op, "mod_4146");
    PMU_IFC mod_4147_bufferize <- mkPMU(2);
    Operation_IFC mod_4147_inner = mod_4147_bufferize.operation;
    Operation_IFC mod_4147 <- mkDebugOperation(mod_4147_inner, "mod_4147");
    Broadcast_IFC#(2) mod_4148_inner <- mkBroadcast(2);
    Operation_IFC mod_4148 <- mkDebugOperation(mod_4148_inner.op, "mod_4148");
    PMU_IFC mod_4149_bufferize <- mkPMU(1);
    Operation_IFC mod_4149_inner = mod_4149_bufferize.operation;
    Operation_IFC mod_4149 <- mkDebugOperation(mod_4149_inner, "mod_4149");
    Operation_IFC mod_4150_inner <- mkBinaryMap(1055, matmul_t_tile);
    Operation_IFC mod_4150 <- mkDebugOperation(mod_4150_inner, "mod_4150");
    Operation_IFC mod_4151_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4151 <- mkDebugOperation(mod_4151_inner, "mod_4151");
    Operation_IFC mod_4152_inner <- mkBinaryMap(1823, mul_tile);
    Operation_IFC mod_4152 <- mkDebugOperation(mod_4152_inner, "mod_4152");
    PMU_IFC mod_4153_bufferize <- mkPMU(1);
    Operation_IFC mod_4153_inner = mod_4153_bufferize.operation;
    Operation_IFC mod_4153 <- mkDebugOperation(mod_4153_inner, "mod_4153");
    Operation_IFC mod_4154_inner <- mkBinaryMap(2361, matmul_t_tile);
    Operation_IFC mod_4154 <- mkDebugOperation(mod_4154_inner, "mod_4154");
    Operation_IFC mod_4155_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4155 <- mkDebugOperation(mod_4155_inner, "mod_4155");
    Operation_IFC mod_4156_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4156 <- mkDebugOperation(mod_4156_inner, "mod_4156");
    Operation_IFC mod_4157_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4157 <- mkDebugOperation(mod_4157_inner, "mod_4157");
    Operation_IFC mod_4158_inner <- mkBinaryMap(2722, mul_tile);
    Operation_IFC mod_4158 <- mkDebugOperation(mod_4158_inner, "mod_4158");
    PMU_IFC mod_4159_bufferize <- mkPMU(1);
    Operation_IFC mod_4159_inner = mod_4159_bufferize.operation;
    Operation_IFC mod_4159 <- mkDebugOperation(mod_4159_inner, "mod_4159");
    PMU_IFC mod_4160_bufferize <- mkPMU(2);
    Operation_IFC mod_4160_inner = mod_4160_bufferize.operation;
    Operation_IFC mod_4160 <- mkDebugOperation(mod_4160_inner, "mod_4160");
    PMU_IFC mod_4161_bufferize <- mkPMU(2);
    Operation_IFC mod_4161_inner = mod_4161_bufferize.operation;
    Operation_IFC mod_4161 <- mkDebugOperation(mod_4161_inner, "mod_4161");
    Operation_IFC mod_4162_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4162 <- mkDebugOperation(mod_4162_inner, "mod_4162");
    Operation_IFC mod_4163_inner <- mkFlatten(1);
    Operation_IFC mod_4163 <- mkDebugOperation(mod_4163_inner, "mod_4163");
    Operation_IFC mod_4164_inner <- mkFlatten(0);
    Operation_IFC mod_4164 <- mkDebugOperation(mod_4164_inner, "mod_4164");
    Operation_IFC mod_4165_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4165 <- mkDebugOperation(mod_4165_inner, "mod_4165");
    Operation_IFC mod_4166_inner <- mkUnaryMap(1695, silu_tile);
    Operation_IFC mod_4166 <- mkDebugOperation(mod_4166_inner, "mod_4166");
    Operation_IFC mod_4167_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4167 <- mkDebugOperation(mod_4167_inner, "mod_4167");
    Operation_IFC mod_4168_inner <- mkBinaryMap(1567, matmul_t_tile);
    Operation_IFC mod_4168 <- mkDebugOperation(mod_4168_inner, "mod_4168");
    PMU_IFC mod_4169_bufferize <- mkPMU(2);
    Operation_IFC mod_4169_inner = mod_4169_bufferize.operation;
    Operation_IFC mod_4169 <- mkDebugOperation(mod_4169_inner, "mod_4169");
    Operation_IFC mod_4170_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4170 <- mkDebugOperation(mod_4170_inner, "mod_4170");
    Operation_IFC mod_4171_inner <- mkFlatten(1);
    Operation_IFC mod_4171 <- mkDebugOperation(mod_4171_inner, "mod_4171");
    Operation_IFC mod_4172_inner <- mkFlatten(0);
    Operation_IFC mod_4172 <- mkDebugOperation(mod_4172_inner, "mod_4172");
    PMU_IFC mod_4173_bufferize <- mkPMU(1);
    Operation_IFC mod_4173_inner = mod_4173_bufferize.operation;
    Operation_IFC mod_4173 <- mkDebugOperation(mod_4173_inner, "mod_4173");
    Operation_IFC mod_4174_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4174 <- mkDebugOperation(mod_4174_inner, "mod_4174");
    PMU_IFC mod_4175_bufferize <- mkPMU(2);
    Operation_IFC mod_4175_inner = mod_4175_bufferize.operation;
    Operation_IFC mod_4175 <- mkDebugOperation(mod_4175_inner, "mod_4175");
    Operation_IFC mod_4176_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4176 <- mkDebugOperation(mod_4176_inner, "mod_4176");
    Operation_IFC mod_4177_inner <- mkFlatten(1);
    Operation_IFC mod_4177 <- mkDebugOperation(mod_4177_inner, "mod_4177");
    Operation_IFC mod_4178_inner <- mkFlatten(0);
    Operation_IFC mod_4178 <- mkDebugOperation(mod_4178_inner, "mod_4178");
    Operation_IFC mod_4179_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4179 <- mkDebugOperation(mod_4179_inner, "mod_4179");
    Operation_IFC mod_4180_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4180 <- mkDebugOperation(mod_4180_inner, "mod_4180");
    PMU_IFC mod_4181_bufferize <- mkPMU(2);
    Operation_IFC mod_4181_inner = mod_4181_bufferize.operation;
    Operation_IFC mod_4181 <- mkDebugOperation(mod_4181_inner, "mod_4181");
    rule rule_5354;
        ChannelMessage t;
        t <- mod_4160.get(0);
        mod_4160.put(1, t);
    endrule
    rule rule_5355;
        ChannelMessage t;
        t <- mod_4159.get(0);
        mod_4159.put(1, t);
    endrule
    rule rule_5356;
        ChannelMessage t;
        t <- mod_4166.get(0);
        mod_4152.put(1, t);
    endrule
    rule rule_5357;
        ChannelMessage t;
        t <- mod_4150.get(0);
        mod_4151.put(0, t);
    endrule
    rule rule_5358;
        ChannelMessage t;
        t <- mod_4153.get(1);
        mod_4154.put(0, t);
    endrule
    rule rule_5359;
        ChannelMessage t;
        t <- mod_4161.get(1);
        mod_4154.put(1, t);
    endrule
    rule rule_5360;
        ChannelMessage t;
        t <- mod_4178.get(0);
        mod_4177.put(0, t);
    endrule
    rule rule_5361;
        ChannelMessage t;
        t <- mod_4164.get(0);
        mod_4163.put(0, t);
    endrule
    rule rule_5362;
        ChannelMessage t;
        t <- mod_4143.get(0);
        mod_4144.put(0, t);
    endrule
    rule rule_5363;
        ChannelMessage t;
        t <- mod_4170.get(0);
        mod_4169.put(1, t);
    endrule
    rule rule_5364;
        ChannelMessage t;
        t <- mod_4151.get(0);
        mod_4152.put(0, t);
    endrule
    rule rule_5365;
        ChannelMessage t;
        t <- mod_4152.get(0);
        mod_4153.put(0, t);
    endrule
    rule rule_5366;
        ChannelMessage t;
        t <- mod_4159.get(1);
        mod_4157.put(1, t);
    endrule
    rule rule_5367;
        ChannelMessage t;
        t <- mod_4157.get(1);
        mod_4158.put(1, t);
    endrule
    rule rule_5368;
        ChannelMessage t;
        t <- mod_4161.get(0);
        mod_4162.put(0, t);
    endrule
    rule rule_5369;
        ChannelMessage t;
        t <- mod_4169.get(0);
        mod_4170.put(0, t);
    endrule
    rule rule_5370;
        ChannelMessage t;
        t <- mod_4174.get(0);
        mod_4173.put(1, t);
    endrule
    rule rule_5371;
        ChannelMessage t;
        t <- mod_4177.get(0);
        mod_4175.put(0, t);
    endrule
    rule rule_5372;
        ChannelMessage t;
        t <- mod_4149.get(0);
        mod_4179.put(0, t);
    endrule
    rule rule_5373;
        ChannelMessage t;
        t <- mod_4142.get(0);
        mod_4143.put(0, t);
    endrule
    rule rule_5374;
        ChannelMessage t;
        t <- mod_4147.get(1);
        mod_4148.put(0, t);
    endrule
    rule rule_5375;
        ChannelMessage t;
        t <- mod_4168.get(0);
        mod_4167.put(0, t);
    endrule
    rule rule_5376;
        ChannelMessage t;
        t <- mod_4156.get(0);
        mod_4160.put(0, t);
    endrule
    rule rule_5377;
        ChannelMessage t;
        t <- mod_4155.get(0);
        mod_4156.put(0, t);
    endrule
    rule rule_5378;
        ChannelMessage t;
        t <- mod_4147.get(0);
        mod_4180.put(0, t);
    endrule
    rule rule_5379;
        ChannelMessage t;
        t <- mod_4148.get(0);
        mod_4173.put(0, t);
    endrule
    rule rule_5380;
        ChannelMessage t;
        t <- mod_4169.get(1);
        mod_4168.put(1, t);
    endrule
    rule rule_5381;
        ChannelMessage t;
        t <- mod_4149.get(1);
        mod_4150.put(0, t);
    endrule
    rule rule_5382;
        ChannelMessage t;
        t <- mod_4154.get(0);
        mod_4155.put(0, t);
    endrule
    rule rule_5383;
        ChannelMessage t;
        t <- mod_4153.get(0);
        mod_4165.put(0, t);
    endrule
    rule rule_5384;
        ChannelMessage t;
        t <- mod_4175.get(1);
        mod_4150.put(1, t);
    endrule
    rule rule_5385;
        ChannelMessage t;
        t <- mod_4144.get(0);
        mod_4145.put(0, t);
    endrule
    rule rule_5386;
        ChannelMessage t;
        t <- mod_4167.get(0);
        mod_4166.put(0, t);
    endrule
    rule rule_5387;
        ChannelMessage t;
        t <- mod_4163.get(0);
        mod_4161.put(0, t);
    endrule
    rule rule_5388;
        ChannelMessage t;
        t <- mod_4145.get(1);
        mod_4146.put(0, t);
    endrule
    rule rule_5389;
        ChannelMessage t;
        t <- mod_4175.get(0);
        mod_4176.put(0, t);
    endrule
    rule rule_5390;
        ChannelMessage t;
        t <- mod_4173.get(0);
        mod_4174.put(0, t);
    endrule
    rule rule_5391;
        ChannelMessage t;
        t <- mod_4171.get(0);
        mod_4169.put(0, t);
    endrule
    rule rule_5392;
        ChannelMessage t;
        t <- mod_4181.get(1);
        mod_4145.put(1, t);
    endrule
    rule rule_5393;
        ChannelMessage t;
        t <- mod_4148.get(1);
        mod_4149.put(0, t);
    endrule
    rule rule_5394;
        ChannelMessage t;
        t <- mod_4157.get(0);
        mod_4159.put(0, t);
    endrule
    rule rule_5395;
        ChannelMessage t;
        t <- mod_4146.get(3);
        mod_4147.put(0, t);
    endrule
    rule rule_5396;
        ChannelMessage t;
        t <- mod_4145.get(0);
        mod_4181.put(0, t);
    endrule
    rule rule_5397;
        ChannelMessage t;
        t <- mod_4179.get(0);
        mod_4149.put(1, t);
    endrule
    rule rule_5398;
        ChannelMessage t;
        t <- mod_4176.get(0);
        mod_4175.put(1, t);
    endrule
    rule rule_5399;
        ChannelMessage t;
        t <- mod_4160.get(1);
        mod_4156.put(1, t);
    endrule
    rule rule_5400;
        ChannelMessage t;
        t <- mod_4165.get(0);
        mod_4153.put(1, t);
    endrule
    rule rule_5401;
        ChannelMessage t;
        t <- mod_4156.get(1);
        mod_4157.put(0, t);
    endrule
    rule rule_5402;
        ChannelMessage t;
        t <- mod_4162.get(0);
        mod_4161.put(1, t);
    endrule
    rule rule_5403;
        ChannelMessage t;
        t <- mod_4181.get(0);
        mod_4181.put(1, t);
    endrule
    rule rule_5404;
        ChannelMessage t;
        t <- mod_4180.get(0);
        mod_4147.put(1, t);
    endrule
    rule rule_5405;
        ChannelMessage t;
        t <- mod_4173.get(1);
        mod_4168.put(0, t);
    endrule
    rule rule_5406;
        ChannelMessage t;
        t <- mod_4172.get(0);
        mod_4171.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4142.put(0, t);
        end
        if (i == 1) begin
            mod_4158.put(0, t);
        end
        if (i == 2) begin
            mod_4164.put(0, t);
        end
        if (i == 3) begin
            mod_4172.put(0, t);
        end
        if (i == 4) begin
            mod_4178.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_4146.get(0);
        end
        if (i == 2) begin
            t <- mod_4146.get(1);
        end
        if (i == 3) begin
            t <- mod_4146.get(2);
        end
        if (i == 1) begin
            t <- mod_4158.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6136 (Operation_IFC);
    Operation_IFC mod_4183_inner <- mkReshape(2, 64);
    Operation_IFC mod_4183 <- mkDebugOperation(mod_4183_inner, "mod_4183");
    Operation_IFC mod_4184_inner <- mkFlatten(1);
    Operation_IFC mod_4184 <- mkDebugOperation(mod_4184_inner, "mod_4184");
    Operation_IFC mod_4185_inner <- mkFlatten(2);
    Operation_IFC mod_4185 <- mkDebugOperation(mod_4185_inner, "mod_4185");
    Operation_IFC mod_4186_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4186 <- mkDebugOperation(mod_4186_inner, "mod_4186");
    Broadcast_IFC#(4) mod_4187_inner <- mkBroadcast(4);
    Operation_IFC mod_4187 <- mkDebugOperation(mod_4187_inner.op, "mod_4187");
    PMU_IFC mod_4188_bufferize <- mkPMU(2);
    Operation_IFC mod_4188_inner = mod_4188_bufferize.operation;
    Operation_IFC mod_4188 <- mkDebugOperation(mod_4188_inner, "mod_4188");
    Broadcast_IFC#(2) mod_4189_inner <- mkBroadcast(2);
    Operation_IFC mod_4189 <- mkDebugOperation(mod_4189_inner.op, "mod_4189");
    PMU_IFC mod_4190_bufferize <- mkPMU(1);
    Operation_IFC mod_4190_inner = mod_4190_bufferize.operation;
    Operation_IFC mod_4190 <- mkDebugOperation(mod_4190_inner, "mod_4190");
    Operation_IFC mod_4191_inner <- mkBinaryMap(1054, matmul_t_tile);
    Operation_IFC mod_4191 <- mkDebugOperation(mod_4191_inner, "mod_4191");
    Operation_IFC mod_4192_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4192 <- mkDebugOperation(mod_4192_inner, "mod_4192");
    Operation_IFC mod_4193_inner <- mkBinaryMap(1822, mul_tile);
    Operation_IFC mod_4193 <- mkDebugOperation(mod_4193_inner, "mod_4193");
    PMU_IFC mod_4194_bufferize <- mkPMU(1);
    Operation_IFC mod_4194_inner = mod_4194_bufferize.operation;
    Operation_IFC mod_4194 <- mkDebugOperation(mod_4194_inner, "mod_4194");
    Operation_IFC mod_4195_inner <- mkBinaryMap(2359, matmul_t_tile);
    Operation_IFC mod_4195 <- mkDebugOperation(mod_4195_inner, "mod_4195");
    Operation_IFC mod_4196_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4196 <- mkDebugOperation(mod_4196_inner, "mod_4196");
    Operation_IFC mod_4197_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4197 <- mkDebugOperation(mod_4197_inner, "mod_4197");
    Operation_IFC mod_4198_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4198 <- mkDebugOperation(mod_4198_inner, "mod_4198");
    Operation_IFC mod_4199_inner <- mkBinaryMap(2721, mul_tile);
    Operation_IFC mod_4199 <- mkDebugOperation(mod_4199_inner, "mod_4199");
    PMU_IFC mod_4200_bufferize <- mkPMU(1);
    Operation_IFC mod_4200_inner = mod_4200_bufferize.operation;
    Operation_IFC mod_4200 <- mkDebugOperation(mod_4200_inner, "mod_4200");
    PMU_IFC mod_4201_bufferize <- mkPMU(2);
    Operation_IFC mod_4201_inner = mod_4201_bufferize.operation;
    Operation_IFC mod_4201 <- mkDebugOperation(mod_4201_inner, "mod_4201");
    PMU_IFC mod_4202_bufferize <- mkPMU(2);
    Operation_IFC mod_4202_inner = mod_4202_bufferize.operation;
    Operation_IFC mod_4202 <- mkDebugOperation(mod_4202_inner, "mod_4202");
    Operation_IFC mod_4203_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4203 <- mkDebugOperation(mod_4203_inner, "mod_4203");
    Operation_IFC mod_4204_inner <- mkFlatten(1);
    Operation_IFC mod_4204 <- mkDebugOperation(mod_4204_inner, "mod_4204");
    Operation_IFC mod_4205_inner <- mkFlatten(0);
    Operation_IFC mod_4205 <- mkDebugOperation(mod_4205_inner, "mod_4205");
    Operation_IFC mod_4206_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4206 <- mkDebugOperation(mod_4206_inner, "mod_4206");
    Operation_IFC mod_4207_inner <- mkUnaryMap(1694, silu_tile);
    Operation_IFC mod_4207 <- mkDebugOperation(mod_4207_inner, "mod_4207");
    Operation_IFC mod_4208_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4208 <- mkDebugOperation(mod_4208_inner, "mod_4208");
    Operation_IFC mod_4209_inner <- mkBinaryMap(1566, matmul_t_tile);
    Operation_IFC mod_4209 <- mkDebugOperation(mod_4209_inner, "mod_4209");
    PMU_IFC mod_4210_bufferize <- mkPMU(2);
    Operation_IFC mod_4210_inner = mod_4210_bufferize.operation;
    Operation_IFC mod_4210 <- mkDebugOperation(mod_4210_inner, "mod_4210");
    Operation_IFC mod_4211_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4211 <- mkDebugOperation(mod_4211_inner, "mod_4211");
    Operation_IFC mod_4212_inner <- mkFlatten(1);
    Operation_IFC mod_4212 <- mkDebugOperation(mod_4212_inner, "mod_4212");
    Operation_IFC mod_4213_inner <- mkFlatten(0);
    Operation_IFC mod_4213 <- mkDebugOperation(mod_4213_inner, "mod_4213");
    PMU_IFC mod_4214_bufferize <- mkPMU(1);
    Operation_IFC mod_4214_inner = mod_4214_bufferize.operation;
    Operation_IFC mod_4214 <- mkDebugOperation(mod_4214_inner, "mod_4214");
    Operation_IFC mod_4215_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4215 <- mkDebugOperation(mod_4215_inner, "mod_4215");
    PMU_IFC mod_4216_bufferize <- mkPMU(2);
    Operation_IFC mod_4216_inner = mod_4216_bufferize.operation;
    Operation_IFC mod_4216 <- mkDebugOperation(mod_4216_inner, "mod_4216");
    Operation_IFC mod_4217_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4217 <- mkDebugOperation(mod_4217_inner, "mod_4217");
    Operation_IFC mod_4218_inner <- mkFlatten(1);
    Operation_IFC mod_4218 <- mkDebugOperation(mod_4218_inner, "mod_4218");
    Operation_IFC mod_4219_inner <- mkFlatten(0);
    Operation_IFC mod_4219 <- mkDebugOperation(mod_4219_inner, "mod_4219");
    Operation_IFC mod_4220_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4220 <- mkDebugOperation(mod_4220_inner, "mod_4220");
    Operation_IFC mod_4221_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4221 <- mkDebugOperation(mod_4221_inner, "mod_4221");
    PMU_IFC mod_4222_bufferize <- mkPMU(2);
    Operation_IFC mod_4222_inner = mod_4222_bufferize.operation;
    Operation_IFC mod_4222 <- mkDebugOperation(mod_4222_inner, "mod_4222");
    rule rule_5407;
        ChannelMessage t;
        t <- mod_4186.get(1);
        mod_4187.put(0, t);
    endrule
    rule rule_5408;
        ChannelMessage t;
        t <- mod_4197.get(0);
        mod_4201.put(0, t);
    endrule
    rule rule_5409;
        ChannelMessage t;
        t <- mod_4187.get(3);
        mod_4188.put(0, t);
    endrule
    rule rule_5410;
        ChannelMessage t;
        t <- mod_4221.get(0);
        mod_4188.put(1, t);
    endrule
    rule rule_5411;
        ChannelMessage t;
        t <- mod_4201.get(1);
        mod_4197.put(1, t);
    endrule
    rule rule_5412;
        ChannelMessage t;
        t <- mod_4202.get(0);
        mod_4203.put(0, t);
    endrule
    rule rule_5413;
        ChannelMessage t;
        t <- mod_4204.get(0);
        mod_4202.put(0, t);
    endrule
    rule rule_5414;
        ChannelMessage t;
        t <- mod_4188.get(0);
        mod_4221.put(0, t);
    endrule
    rule rule_5415;
        ChannelMessage t;
        t <- mod_4212.get(0);
        mod_4210.put(0, t);
    endrule
    rule rule_5416;
        ChannelMessage t;
        t <- mod_4184.get(0);
        mod_4185.put(0, t);
    endrule
    rule rule_5417;
        ChannelMessage t;
        t <- mod_4188.get(1);
        mod_4189.put(0, t);
    endrule
    rule rule_5418;
        ChannelMessage t;
        t <- mod_4189.get(0);
        mod_4214.put(0, t);
    endrule
    rule rule_5419;
        ChannelMessage t;
        t <- mod_4202.get(1);
        mod_4195.put(1, t);
    endrule
    rule rule_5420;
        ChannelMessage t;
        t <- mod_4218.get(0);
        mod_4216.put(0, t);
    endrule
    rule rule_5421;
        ChannelMessage t;
        t <- mod_4190.get(0);
        mod_4220.put(0, t);
    endrule
    rule rule_5422;
        ChannelMessage t;
        t <- mod_4214.get(0);
        mod_4215.put(0, t);
    endrule
    rule rule_5423;
        ChannelMessage t;
        t <- mod_4198.get(1);
        mod_4199.put(1, t);
    endrule
    rule rule_5424;
        ChannelMessage t;
        t <- mod_4191.get(0);
        mod_4192.put(0, t);
    endrule
    rule rule_5425;
        ChannelMessage t;
        t <- mod_4194.get(0);
        mod_4206.put(0, t);
    endrule
    rule rule_5426;
        ChannelMessage t;
        t <- mod_4190.get(1);
        mod_4191.put(0, t);
    endrule
    rule rule_5427;
        ChannelMessage t;
        t <- mod_4194.get(1);
        mod_4195.put(0, t);
    endrule
    rule rule_5428;
        ChannelMessage t;
        t <- mod_4207.get(0);
        mod_4193.put(1, t);
    endrule
    rule rule_5429;
        ChannelMessage t;
        t <- mod_4205.get(0);
        mod_4204.put(0, t);
    endrule
    rule rule_5430;
        ChannelMessage t;
        t <- mod_4208.get(0);
        mod_4207.put(0, t);
    endrule
    rule rule_5431;
        ChannelMessage t;
        t <- mod_4185.get(0);
        mod_4186.put(0, t);
    endrule
    rule rule_5432;
        ChannelMessage t;
        t <- mod_4206.get(0);
        mod_4194.put(1, t);
    endrule
    rule rule_5433;
        ChannelMessage t;
        t <- mod_4213.get(0);
        mod_4212.put(0, t);
    endrule
    rule rule_5434;
        ChannelMessage t;
        t <- mod_4222.get(1);
        mod_4186.put(1, t);
    endrule
    rule rule_5435;
        ChannelMessage t;
        t <- mod_4189.get(1);
        mod_4190.put(0, t);
    endrule
    rule rule_5436;
        ChannelMessage t;
        t <- mod_4198.get(0);
        mod_4200.put(0, t);
    endrule
    rule rule_5437;
        ChannelMessage t;
        t <- mod_4215.get(0);
        mod_4214.put(1, t);
    endrule
    rule rule_5438;
        ChannelMessage t;
        t <- mod_4193.get(0);
        mod_4194.put(0, t);
    endrule
    rule rule_5439;
        ChannelMessage t;
        t <- mod_4210.get(0);
        mod_4211.put(0, t);
    endrule
    rule rule_5440;
        ChannelMessage t;
        t <- mod_4200.get(1);
        mod_4198.put(1, t);
    endrule
    rule rule_5441;
        ChannelMessage t;
        t <- mod_4197.get(1);
        mod_4198.put(0, t);
    endrule
    rule rule_5442;
        ChannelMessage t;
        t <- mod_4200.get(0);
        mod_4200.put(1, t);
    endrule
    rule rule_5443;
        ChannelMessage t;
        t <- mod_4201.get(0);
        mod_4201.put(1, t);
    endrule
    rule rule_5444;
        ChannelMessage t;
        t <- mod_4211.get(0);
        mod_4210.put(1, t);
    endrule
    rule rule_5445;
        ChannelMessage t;
        t <- mod_4220.get(0);
        mod_4190.put(1, t);
    endrule
    rule rule_5446;
        ChannelMessage t;
        t <- mod_4214.get(1);
        mod_4209.put(0, t);
    endrule
    rule rule_5447;
        ChannelMessage t;
        t <- mod_4196.get(0);
        mod_4197.put(0, t);
    endrule
    rule rule_5448;
        ChannelMessage t;
        t <- mod_4209.get(0);
        mod_4208.put(0, t);
    endrule
    rule rule_5449;
        ChannelMessage t;
        t <- mod_4222.get(0);
        mod_4222.put(1, t);
    endrule
    rule rule_5450;
        ChannelMessage t;
        t <- mod_4216.get(1);
        mod_4191.put(1, t);
    endrule
    rule rule_5451;
        ChannelMessage t;
        t <- mod_4186.get(0);
        mod_4222.put(0, t);
    endrule
    rule rule_5452;
        ChannelMessage t;
        t <- mod_4183.get(0);
        mod_4184.put(0, t);
    endrule
    rule rule_5453;
        ChannelMessage t;
        t <- mod_4192.get(0);
        mod_4193.put(0, t);
    endrule
    rule rule_5454;
        ChannelMessage t;
        t <- mod_4210.get(1);
        mod_4209.put(1, t);
    endrule
    rule rule_5455;
        ChannelMessage t;
        t <- mod_4216.get(0);
        mod_4217.put(0, t);
    endrule
    rule rule_5456;
        ChannelMessage t;
        t <- mod_4195.get(0);
        mod_4196.put(0, t);
    endrule
    rule rule_5457;
        ChannelMessage t;
        t <- mod_4203.get(0);
        mod_4202.put(1, t);
    endrule
    rule rule_5458;
        ChannelMessage t;
        t <- mod_4217.get(0);
        mod_4216.put(1, t);
    endrule
    rule rule_5459;
        ChannelMessage t;
        t <- mod_4219.get(0);
        mod_4218.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4183.put(0, t);
        end
        if (i == 1) begin
            mod_4199.put(0, t);
        end
        if (i == 2) begin
            mod_4205.put(0, t);
        end
        if (i == 3) begin
            mod_4213.put(0, t);
        end
        if (i == 4) begin
            mod_4219.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_4187.get(0);
        end
        if (i == 1) begin
            t <- mod_4187.get(1);
        end
        if (i == 2) begin
            t <- mod_4187.get(2);
        end
        if (i == 3) begin
            t <- mod_4199.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6137 (Operation_IFC);
    Operation_IFC mod_4224_inner <- mkReshape(2, 64);
    Operation_IFC mod_4224 <- mkDebugOperation(mod_4224_inner, "mod_4224");
    Operation_IFC mod_4225_inner <- mkFlatten(1);
    Operation_IFC mod_4225 <- mkDebugOperation(mod_4225_inner, "mod_4225");
    Operation_IFC mod_4226_inner <- mkFlatten(2);
    Operation_IFC mod_4226 <- mkDebugOperation(mod_4226_inner, "mod_4226");
    Operation_IFC mod_4227_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4227 <- mkDebugOperation(mod_4227_inner, "mod_4227");
    Broadcast_IFC#(4) mod_4228_inner <- mkBroadcast(4);
    Operation_IFC mod_4228 <- mkDebugOperation(mod_4228_inner.op, "mod_4228");
    PMU_IFC mod_4229_bufferize <- mkPMU(2);
    Operation_IFC mod_4229_inner = mod_4229_bufferize.operation;
    Operation_IFC mod_4229 <- mkDebugOperation(mod_4229_inner, "mod_4229");
    Broadcast_IFC#(2) mod_4230_inner <- mkBroadcast(2);
    Operation_IFC mod_4230 <- mkDebugOperation(mod_4230_inner.op, "mod_4230");
    PMU_IFC mod_4231_bufferize <- mkPMU(1);
    Operation_IFC mod_4231_inner = mod_4231_bufferize.operation;
    Operation_IFC mod_4231 <- mkDebugOperation(mod_4231_inner, "mod_4231");
    Operation_IFC mod_4232_inner <- mkBinaryMap(1053, matmul_t_tile);
    Operation_IFC mod_4232 <- mkDebugOperation(mod_4232_inner, "mod_4232");
    Operation_IFC mod_4233_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4233 <- mkDebugOperation(mod_4233_inner, "mod_4233");
    Operation_IFC mod_4234_inner <- mkBinaryMap(1821, mul_tile);
    Operation_IFC mod_4234 <- mkDebugOperation(mod_4234_inner, "mod_4234");
    PMU_IFC mod_4235_bufferize <- mkPMU(1);
    Operation_IFC mod_4235_inner = mod_4235_bufferize.operation;
    Operation_IFC mod_4235 <- mkDebugOperation(mod_4235_inner, "mod_4235");
    Operation_IFC mod_4236_inner <- mkBinaryMap(2357, matmul_t_tile);
    Operation_IFC mod_4236 <- mkDebugOperation(mod_4236_inner, "mod_4236");
    Operation_IFC mod_4237_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4237 <- mkDebugOperation(mod_4237_inner, "mod_4237");
    Operation_IFC mod_4238_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4238 <- mkDebugOperation(mod_4238_inner, "mod_4238");
    Operation_IFC mod_4239_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4239 <- mkDebugOperation(mod_4239_inner, "mod_4239");
    Operation_IFC mod_4240_inner <- mkBinaryMap(2720, mul_tile);
    Operation_IFC mod_4240 <- mkDebugOperation(mod_4240_inner, "mod_4240");
    PMU_IFC mod_4241_bufferize <- mkPMU(1);
    Operation_IFC mod_4241_inner = mod_4241_bufferize.operation;
    Operation_IFC mod_4241 <- mkDebugOperation(mod_4241_inner, "mod_4241");
    PMU_IFC mod_4242_bufferize <- mkPMU(2);
    Operation_IFC mod_4242_inner = mod_4242_bufferize.operation;
    Operation_IFC mod_4242 <- mkDebugOperation(mod_4242_inner, "mod_4242");
    PMU_IFC mod_4243_bufferize <- mkPMU(2);
    Operation_IFC mod_4243_inner = mod_4243_bufferize.operation;
    Operation_IFC mod_4243 <- mkDebugOperation(mod_4243_inner, "mod_4243");
    Operation_IFC mod_4244_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4244 <- mkDebugOperation(mod_4244_inner, "mod_4244");
    Operation_IFC mod_4245_inner <- mkFlatten(1);
    Operation_IFC mod_4245 <- mkDebugOperation(mod_4245_inner, "mod_4245");
    Operation_IFC mod_4246_inner <- mkFlatten(0);
    Operation_IFC mod_4246 <- mkDebugOperation(mod_4246_inner, "mod_4246");
    Operation_IFC mod_4247_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4247 <- mkDebugOperation(mod_4247_inner, "mod_4247");
    Operation_IFC mod_4248_inner <- mkUnaryMap(1693, silu_tile);
    Operation_IFC mod_4248 <- mkDebugOperation(mod_4248_inner, "mod_4248");
    Operation_IFC mod_4249_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4249 <- mkDebugOperation(mod_4249_inner, "mod_4249");
    Operation_IFC mod_4250_inner <- mkBinaryMap(1565, matmul_t_tile);
    Operation_IFC mod_4250 <- mkDebugOperation(mod_4250_inner, "mod_4250");
    PMU_IFC mod_4251_bufferize <- mkPMU(2);
    Operation_IFC mod_4251_inner = mod_4251_bufferize.operation;
    Operation_IFC mod_4251 <- mkDebugOperation(mod_4251_inner, "mod_4251");
    Operation_IFC mod_4252_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4252 <- mkDebugOperation(mod_4252_inner, "mod_4252");
    Operation_IFC mod_4253_inner <- mkFlatten(1);
    Operation_IFC mod_4253 <- mkDebugOperation(mod_4253_inner, "mod_4253");
    Operation_IFC mod_4254_inner <- mkFlatten(0);
    Operation_IFC mod_4254 <- mkDebugOperation(mod_4254_inner, "mod_4254");
    PMU_IFC mod_4255_bufferize <- mkPMU(1);
    Operation_IFC mod_4255_inner = mod_4255_bufferize.operation;
    Operation_IFC mod_4255 <- mkDebugOperation(mod_4255_inner, "mod_4255");
    Operation_IFC mod_4256_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4256 <- mkDebugOperation(mod_4256_inner, "mod_4256");
    PMU_IFC mod_4257_bufferize <- mkPMU(2);
    Operation_IFC mod_4257_inner = mod_4257_bufferize.operation;
    Operation_IFC mod_4257 <- mkDebugOperation(mod_4257_inner, "mod_4257");
    Operation_IFC mod_4258_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4258 <- mkDebugOperation(mod_4258_inner, "mod_4258");
    Operation_IFC mod_4259_inner <- mkFlatten(1);
    Operation_IFC mod_4259 <- mkDebugOperation(mod_4259_inner, "mod_4259");
    Operation_IFC mod_4260_inner <- mkFlatten(0);
    Operation_IFC mod_4260 <- mkDebugOperation(mod_4260_inner, "mod_4260");
    Operation_IFC mod_4261_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4261 <- mkDebugOperation(mod_4261_inner, "mod_4261");
    Operation_IFC mod_4262_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4262 <- mkDebugOperation(mod_4262_inner, "mod_4262");
    PMU_IFC mod_4263_bufferize <- mkPMU(2);
    Operation_IFC mod_4263_inner = mod_4263_bufferize.operation;
    Operation_IFC mod_4263 <- mkDebugOperation(mod_4263_inner, "mod_4263");
    rule rule_5460;
        ChannelMessage t;
        t <- mod_4226.get(0);
        mod_4227.put(0, t);
    endrule
    rule rule_5461;
        ChannelMessage t;
        t <- mod_4250.get(0);
        mod_4249.put(0, t);
    endrule
    rule rule_5462;
        ChannelMessage t;
        t <- mod_4231.get(1);
        mod_4232.put(0, t);
    endrule
    rule rule_5463;
        ChannelMessage t;
        t <- mod_4225.get(0);
        mod_4226.put(0, t);
    endrule
    rule rule_5464;
        ChannelMessage t;
        t <- mod_4230.get(1);
        mod_4231.put(0, t);
    endrule
    rule rule_5465;
        ChannelMessage t;
        t <- mod_4236.get(0);
        mod_4237.put(0, t);
    endrule
    rule rule_5466;
        ChannelMessage t;
        t <- mod_4227.get(1);
        mod_4228.put(0, t);
    endrule
    rule rule_5467;
        ChannelMessage t;
        t <- mod_4243.get(1);
        mod_4236.put(1, t);
    endrule
    rule rule_5468;
        ChannelMessage t;
        t <- mod_4245.get(0);
        mod_4243.put(0, t);
    endrule
    rule rule_5469;
        ChannelMessage t;
        t <- mod_4246.get(0);
        mod_4245.put(0, t);
    endrule
    rule rule_5470;
        ChannelMessage t;
        t <- mod_4252.get(0);
        mod_4251.put(1, t);
    endrule
    rule rule_5471;
        ChannelMessage t;
        t <- mod_4259.get(0);
        mod_4257.put(0, t);
    endrule
    rule rule_5472;
        ChannelMessage t;
        t <- mod_4242.get(1);
        mod_4238.put(1, t);
    endrule
    rule rule_5473;
        ChannelMessage t;
        t <- mod_4260.get(0);
        mod_4259.put(0, t);
    endrule
    rule rule_5474;
        ChannelMessage t;
        t <- mod_4257.get(1);
        mod_4232.put(1, t);
    endrule
    rule rule_5475;
        ChannelMessage t;
        t <- mod_4235.get(1);
        mod_4236.put(0, t);
    endrule
    rule rule_5476;
        ChannelMessage t;
        t <- mod_4239.get(0);
        mod_4241.put(0, t);
    endrule
    rule rule_5477;
        ChannelMessage t;
        t <- mod_4255.get(0);
        mod_4256.put(0, t);
    endrule
    rule rule_5478;
        ChannelMessage t;
        t <- mod_4247.get(0);
        mod_4235.put(1, t);
    endrule
    rule rule_5479;
        ChannelMessage t;
        t <- mod_4238.get(1);
        mod_4239.put(0, t);
    endrule
    rule rule_5480;
        ChannelMessage t;
        t <- mod_4256.get(0);
        mod_4255.put(1, t);
    endrule
    rule rule_5481;
        ChannelMessage t;
        t <- mod_4237.get(0);
        mod_4238.put(0, t);
    endrule
    rule rule_5482;
        ChannelMessage t;
        t <- mod_4235.get(0);
        mod_4247.put(0, t);
    endrule
    rule rule_5483;
        ChannelMessage t;
        t <- mod_4262.get(0);
        mod_4229.put(1, t);
    endrule
    rule rule_5484;
        ChannelMessage t;
        t <- mod_4229.get(1);
        mod_4230.put(0, t);
    endrule
    rule rule_5485;
        ChannelMessage t;
        t <- mod_4254.get(0);
        mod_4253.put(0, t);
    endrule
    rule rule_5486;
        ChannelMessage t;
        t <- mod_4229.get(0);
        mod_4262.put(0, t);
    endrule
    rule rule_5487;
        ChannelMessage t;
        t <- mod_4227.get(0);
        mod_4263.put(0, t);
    endrule
    rule rule_5488;
        ChannelMessage t;
        t <- mod_4253.get(0);
        mod_4251.put(0, t);
    endrule
    rule rule_5489;
        ChannelMessage t;
        t <- mod_4230.get(0);
        mod_4255.put(0, t);
    endrule
    rule rule_5490;
        ChannelMessage t;
        t <- mod_4257.get(0);
        mod_4258.put(0, t);
    endrule
    rule rule_5491;
        ChannelMessage t;
        t <- mod_4224.get(0);
        mod_4225.put(0, t);
    endrule
    rule rule_5492;
        ChannelMessage t;
        t <- mod_4242.get(0);
        mod_4242.put(1, t);
    endrule
    rule rule_5493;
        ChannelMessage t;
        t <- mod_4234.get(0);
        mod_4235.put(0, t);
    endrule
    rule rule_5494;
        ChannelMessage t;
        t <- mod_4233.get(0);
        mod_4234.put(0, t);
    endrule
    rule rule_5495;
        ChannelMessage t;
        t <- mod_4228.get(3);
        mod_4229.put(0, t);
    endrule
    rule rule_5496;
        ChannelMessage t;
        t <- mod_4232.get(0);
        mod_4233.put(0, t);
    endrule
    rule rule_5497;
        ChannelMessage t;
        t <- mod_4258.get(0);
        mod_4257.put(1, t);
    endrule
    rule rule_5498;
        ChannelMessage t;
        t <- mod_4241.get(1);
        mod_4239.put(1, t);
    endrule
    rule rule_5499;
        ChannelMessage t;
        t <- mod_4231.get(0);
        mod_4261.put(0, t);
    endrule
    rule rule_5500;
        ChannelMessage t;
        t <- mod_4249.get(0);
        mod_4248.put(0, t);
    endrule
    rule rule_5501;
        ChannelMessage t;
        t <- mod_4261.get(0);
        mod_4231.put(1, t);
    endrule
    rule rule_5502;
        ChannelMessage t;
        t <- mod_4241.get(0);
        mod_4241.put(1, t);
    endrule
    rule rule_5503;
        ChannelMessage t;
        t <- mod_4239.get(1);
        mod_4240.put(1, t);
    endrule
    rule rule_5504;
        ChannelMessage t;
        t <- mod_4238.get(0);
        mod_4242.put(0, t);
    endrule
    rule rule_5505;
        ChannelMessage t;
        t <- mod_4255.get(1);
        mod_4250.put(0, t);
    endrule
    rule rule_5506;
        ChannelMessage t;
        t <- mod_4244.get(0);
        mod_4243.put(1, t);
    endrule
    rule rule_5507;
        ChannelMessage t;
        t <- mod_4251.get(1);
        mod_4250.put(1, t);
    endrule
    rule rule_5508;
        ChannelMessage t;
        t <- mod_4243.get(0);
        mod_4244.put(0, t);
    endrule
    rule rule_5509;
        ChannelMessage t;
        t <- mod_4248.get(0);
        mod_4234.put(1, t);
    endrule
    rule rule_5510;
        ChannelMessage t;
        t <- mod_4251.get(0);
        mod_4252.put(0, t);
    endrule
    rule rule_5511;
        ChannelMessage t;
        t <- mod_4263.get(1);
        mod_4227.put(1, t);
    endrule
    rule rule_5512;
        ChannelMessage t;
        t <- mod_4263.get(0);
        mod_4263.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4224.put(0, t);
        end
        if (i == 1) begin
            mod_4240.put(0, t);
        end
        if (i == 2) begin
            mod_4246.put(0, t);
        end
        if (i == 3) begin
            mod_4254.put(0, t);
        end
        if (i == 4) begin
            mod_4260.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_4228.get(0);
        end
        if (i == 3) begin
            t <- mod_4228.get(1);
        end
        if (i == 1) begin
            t <- mod_4228.get(2);
        end
        if (i == 2) begin
            t <- mod_4240.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6138 (Operation_IFC);
    Operation_IFC mod_4265_inner <- mkReshape(2, 64);
    Operation_IFC mod_4265 <- mkDebugOperation(mod_4265_inner, "mod_4265");
    Operation_IFC mod_4266_inner <- mkFlatten(1);
    Operation_IFC mod_4266 <- mkDebugOperation(mod_4266_inner, "mod_4266");
    Operation_IFC mod_4267_inner <- mkFlatten(2);
    Operation_IFC mod_4267 <- mkDebugOperation(mod_4267_inner, "mod_4267");
    Operation_IFC mod_4268_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4268 <- mkDebugOperation(mod_4268_inner, "mod_4268");
    Broadcast_IFC#(4) mod_4269_inner <- mkBroadcast(4);
    Operation_IFC mod_4269 <- mkDebugOperation(mod_4269_inner.op, "mod_4269");
    PMU_IFC mod_4270_bufferize <- mkPMU(2);
    Operation_IFC mod_4270_inner = mod_4270_bufferize.operation;
    Operation_IFC mod_4270 <- mkDebugOperation(mod_4270_inner, "mod_4270");
    Broadcast_IFC#(2) mod_4271_inner <- mkBroadcast(2);
    Operation_IFC mod_4271 <- mkDebugOperation(mod_4271_inner.op, "mod_4271");
    PMU_IFC mod_4272_bufferize <- mkPMU(1);
    Operation_IFC mod_4272_inner = mod_4272_bufferize.operation;
    Operation_IFC mod_4272 <- mkDebugOperation(mod_4272_inner, "mod_4272");
    Operation_IFC mod_4273_inner <- mkBinaryMap(1052, matmul_t_tile);
    Operation_IFC mod_4273 <- mkDebugOperation(mod_4273_inner, "mod_4273");
    Operation_IFC mod_4274_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4274 <- mkDebugOperation(mod_4274_inner, "mod_4274");
    Operation_IFC mod_4275_inner <- mkBinaryMap(1820, mul_tile);
    Operation_IFC mod_4275 <- mkDebugOperation(mod_4275_inner, "mod_4275");
    PMU_IFC mod_4276_bufferize <- mkPMU(1);
    Operation_IFC mod_4276_inner = mod_4276_bufferize.operation;
    Operation_IFC mod_4276 <- mkDebugOperation(mod_4276_inner, "mod_4276");
    Operation_IFC mod_4277_inner <- mkBinaryMap(2355, matmul_t_tile);
    Operation_IFC mod_4277 <- mkDebugOperation(mod_4277_inner, "mod_4277");
    Operation_IFC mod_4278_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4278 <- mkDebugOperation(mod_4278_inner, "mod_4278");
    Operation_IFC mod_4279_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4279 <- mkDebugOperation(mod_4279_inner, "mod_4279");
    Operation_IFC mod_4280_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4280 <- mkDebugOperation(mod_4280_inner, "mod_4280");
    Operation_IFC mod_4281_inner <- mkBinaryMap(2719, mul_tile);
    Operation_IFC mod_4281 <- mkDebugOperation(mod_4281_inner, "mod_4281");
    PMU_IFC mod_4282_bufferize <- mkPMU(1);
    Operation_IFC mod_4282_inner = mod_4282_bufferize.operation;
    Operation_IFC mod_4282 <- mkDebugOperation(mod_4282_inner, "mod_4282");
    PMU_IFC mod_4283_bufferize <- mkPMU(2);
    Operation_IFC mod_4283_inner = mod_4283_bufferize.operation;
    Operation_IFC mod_4283 <- mkDebugOperation(mod_4283_inner, "mod_4283");
    PMU_IFC mod_4284_bufferize <- mkPMU(2);
    Operation_IFC mod_4284_inner = mod_4284_bufferize.operation;
    Operation_IFC mod_4284 <- mkDebugOperation(mod_4284_inner, "mod_4284");
    Operation_IFC mod_4285_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4285 <- mkDebugOperation(mod_4285_inner, "mod_4285");
    Operation_IFC mod_4286_inner <- mkFlatten(1);
    Operation_IFC mod_4286 <- mkDebugOperation(mod_4286_inner, "mod_4286");
    Operation_IFC mod_4287_inner <- mkFlatten(0);
    Operation_IFC mod_4287 <- mkDebugOperation(mod_4287_inner, "mod_4287");
    Operation_IFC mod_4288_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4288 <- mkDebugOperation(mod_4288_inner, "mod_4288");
    Operation_IFC mod_4289_inner <- mkUnaryMap(1692, silu_tile);
    Operation_IFC mod_4289 <- mkDebugOperation(mod_4289_inner, "mod_4289");
    Operation_IFC mod_4290_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4290 <- mkDebugOperation(mod_4290_inner, "mod_4290");
    Operation_IFC mod_4291_inner <- mkBinaryMap(1564, matmul_t_tile);
    Operation_IFC mod_4291 <- mkDebugOperation(mod_4291_inner, "mod_4291");
    PMU_IFC mod_4292_bufferize <- mkPMU(2);
    Operation_IFC mod_4292_inner = mod_4292_bufferize.operation;
    Operation_IFC mod_4292 <- mkDebugOperation(mod_4292_inner, "mod_4292");
    Operation_IFC mod_4293_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4293 <- mkDebugOperation(mod_4293_inner, "mod_4293");
    Operation_IFC mod_4294_inner <- mkFlatten(1);
    Operation_IFC mod_4294 <- mkDebugOperation(mod_4294_inner, "mod_4294");
    Operation_IFC mod_4295_inner <- mkFlatten(0);
    Operation_IFC mod_4295 <- mkDebugOperation(mod_4295_inner, "mod_4295");
    PMU_IFC mod_4296_bufferize <- mkPMU(1);
    Operation_IFC mod_4296_inner = mod_4296_bufferize.operation;
    Operation_IFC mod_4296 <- mkDebugOperation(mod_4296_inner, "mod_4296");
    Operation_IFC mod_4297_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4297 <- mkDebugOperation(mod_4297_inner, "mod_4297");
    PMU_IFC mod_4298_bufferize <- mkPMU(2);
    Operation_IFC mod_4298_inner = mod_4298_bufferize.operation;
    Operation_IFC mod_4298 <- mkDebugOperation(mod_4298_inner, "mod_4298");
    Operation_IFC mod_4299_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4299 <- mkDebugOperation(mod_4299_inner, "mod_4299");
    Operation_IFC mod_4300_inner <- mkFlatten(1);
    Operation_IFC mod_4300 <- mkDebugOperation(mod_4300_inner, "mod_4300");
    Operation_IFC mod_4301_inner <- mkFlatten(0);
    Operation_IFC mod_4301 <- mkDebugOperation(mod_4301_inner, "mod_4301");
    Operation_IFC mod_4302_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4302 <- mkDebugOperation(mod_4302_inner, "mod_4302");
    Operation_IFC mod_4303_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4303 <- mkDebugOperation(mod_4303_inner, "mod_4303");
    PMU_IFC mod_4304_bufferize <- mkPMU(2);
    Operation_IFC mod_4304_inner = mod_4304_bufferize.operation;
    Operation_IFC mod_4304 <- mkDebugOperation(mod_4304_inner, "mod_4304");
    rule rule_5513;
        ChannelMessage t;
        t <- mod_4300.get(0);
        mod_4298.put(0, t);
    endrule
    rule rule_5514;
        ChannelMessage t;
        t <- mod_4280.get(0);
        mod_4282.put(0, t);
    endrule
    rule rule_5515;
        ChannelMessage t;
        t <- mod_4296.get(0);
        mod_4297.put(0, t);
    endrule
    rule rule_5516;
        ChannelMessage t;
        t <- mod_4296.get(1);
        mod_4291.put(0, t);
    endrule
    rule rule_5517;
        ChannelMessage t;
        t <- mod_4273.get(0);
        mod_4274.put(0, t);
    endrule
    rule rule_5518;
        ChannelMessage t;
        t <- mod_4297.get(0);
        mod_4296.put(1, t);
    endrule
    rule rule_5519;
        ChannelMessage t;
        t <- mod_4279.get(0);
        mod_4283.put(0, t);
    endrule
    rule rule_5520;
        ChannelMessage t;
        t <- mod_4285.get(0);
        mod_4284.put(1, t);
    endrule
    rule rule_5521;
        ChannelMessage t;
        t <- mod_4292.get(0);
        mod_4293.put(0, t);
    endrule
    rule rule_5522;
        ChannelMessage t;
        t <- mod_4299.get(0);
        mod_4298.put(1, t);
    endrule
    rule rule_5523;
        ChannelMessage t;
        t <- mod_4268.get(0);
        mod_4304.put(0, t);
    endrule
    rule rule_5524;
        ChannelMessage t;
        t <- mod_4272.get(0);
        mod_4302.put(0, t);
    endrule
    rule rule_5525;
        ChannelMessage t;
        t <- mod_4290.get(0);
        mod_4289.put(0, t);
    endrule
    rule rule_5526;
        ChannelMessage t;
        t <- mod_4298.get(0);
        mod_4299.put(0, t);
    endrule
    rule rule_5527;
        ChannelMessage t;
        t <- mod_4282.get(1);
        mod_4280.put(1, t);
    endrule
    rule rule_5528;
        ChannelMessage t;
        t <- mod_4291.get(0);
        mod_4290.put(0, t);
    endrule
    rule rule_5529;
        ChannelMessage t;
        t <- mod_4282.get(0);
        mod_4282.put(1, t);
    endrule
    rule rule_5530;
        ChannelMessage t;
        t <- mod_4270.get(0);
        mod_4303.put(0, t);
    endrule
    rule rule_5531;
        ChannelMessage t;
        t <- mod_4295.get(0);
        mod_4294.put(0, t);
    endrule
    rule rule_5532;
        ChannelMessage t;
        t <- mod_4304.get(1);
        mod_4268.put(1, t);
    endrule
    rule rule_5533;
        ChannelMessage t;
        t <- mod_4283.get(0);
        mod_4283.put(1, t);
    endrule
    rule rule_5534;
        ChannelMessage t;
        t <- mod_4288.get(0);
        mod_4276.put(1, t);
    endrule
    rule rule_5535;
        ChannelMessage t;
        t <- mod_4304.get(0);
        mod_4304.put(1, t);
    endrule
    rule rule_5536;
        ChannelMessage t;
        t <- mod_4283.get(1);
        mod_4279.put(1, t);
    endrule
    rule rule_5537;
        ChannelMessage t;
        t <- mod_4274.get(0);
        mod_4275.put(0, t);
    endrule
    rule rule_5538;
        ChannelMessage t;
        t <- mod_4275.get(0);
        mod_4276.put(0, t);
    endrule
    rule rule_5539;
        ChannelMessage t;
        t <- mod_4292.get(1);
        mod_4291.put(1, t);
    endrule
    rule rule_5540;
        ChannelMessage t;
        t <- mod_4284.get(0);
        mod_4285.put(0, t);
    endrule
    rule rule_5541;
        ChannelMessage t;
        t <- mod_4267.get(0);
        mod_4268.put(0, t);
    endrule
    rule rule_5542;
        ChannelMessage t;
        t <- mod_4265.get(0);
        mod_4266.put(0, t);
    endrule
    rule rule_5543;
        ChannelMessage t;
        t <- mod_4286.get(0);
        mod_4284.put(0, t);
    endrule
    rule rule_5544;
        ChannelMessage t;
        t <- mod_4279.get(1);
        mod_4280.put(0, t);
    endrule
    rule rule_5545;
        ChannelMessage t;
        t <- mod_4280.get(1);
        mod_4281.put(1, t);
    endrule
    rule rule_5546;
        ChannelMessage t;
        t <- mod_4284.get(1);
        mod_4277.put(1, t);
    endrule
    rule rule_5547;
        ChannelMessage t;
        t <- mod_4294.get(0);
        mod_4292.put(0, t);
    endrule
    rule rule_5548;
        ChannelMessage t;
        t <- mod_4269.get(3);
        mod_4270.put(0, t);
    endrule
    rule rule_5549;
        ChannelMessage t;
        t <- mod_4298.get(1);
        mod_4273.put(1, t);
    endrule
    rule rule_5550;
        ChannelMessage t;
        t <- mod_4303.get(0);
        mod_4270.put(1, t);
    endrule
    rule rule_5551;
        ChannelMessage t;
        t <- mod_4272.get(1);
        mod_4273.put(0, t);
    endrule
    rule rule_5552;
        ChannelMessage t;
        t <- mod_4276.get(0);
        mod_4288.put(0, t);
    endrule
    rule rule_5553;
        ChannelMessage t;
        t <- mod_4287.get(0);
        mod_4286.put(0, t);
    endrule
    rule rule_5554;
        ChannelMessage t;
        t <- mod_4271.get(0);
        mod_4296.put(0, t);
    endrule
    rule rule_5555;
        ChannelMessage t;
        t <- mod_4266.get(0);
        mod_4267.put(0, t);
    endrule
    rule rule_5556;
        ChannelMessage t;
        t <- mod_4289.get(0);
        mod_4275.put(1, t);
    endrule
    rule rule_5557;
        ChannelMessage t;
        t <- mod_4293.get(0);
        mod_4292.put(1, t);
    endrule
    rule rule_5558;
        ChannelMessage t;
        t <- mod_4302.get(0);
        mod_4272.put(1, t);
    endrule
    rule rule_5559;
        ChannelMessage t;
        t <- mod_4271.get(1);
        mod_4272.put(0, t);
    endrule
    rule rule_5560;
        ChannelMessage t;
        t <- mod_4277.get(0);
        mod_4278.put(0, t);
    endrule
    rule rule_5561;
        ChannelMessage t;
        t <- mod_4270.get(1);
        mod_4271.put(0, t);
    endrule
    rule rule_5562;
        ChannelMessage t;
        t <- mod_4278.get(0);
        mod_4279.put(0, t);
    endrule
    rule rule_5563;
        ChannelMessage t;
        t <- mod_4268.get(1);
        mod_4269.put(0, t);
    endrule
    rule rule_5564;
        ChannelMessage t;
        t <- mod_4276.get(1);
        mod_4277.put(0, t);
    endrule
    rule rule_5565;
        ChannelMessage t;
        t <- mod_4301.get(0);
        mod_4300.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4265.put(0, t);
        end
        if (i == 1) begin
            mod_4281.put(0, t);
        end
        if (i == 2) begin
            mod_4287.put(0, t);
        end
        if (i == 3) begin
            mod_4295.put(0, t);
        end
        if (i == 4) begin
            mod_4301.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_4269.get(0);
        end
        if (i == 1) begin
            t <- mod_4269.get(1);
        end
        if (i == 0) begin
            t <- mod_4269.get(2);
        end
        if (i == 2) begin
            t <- mod_4281.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6139 (Operation_IFC);
    Operation_IFC mod_4306_inner <- mkReshape(2, 64);
    Operation_IFC mod_4306 <- mkDebugOperation(mod_4306_inner, "mod_4306");
    Operation_IFC mod_4307_inner <- mkFlatten(1);
    Operation_IFC mod_4307 <- mkDebugOperation(mod_4307_inner, "mod_4307");
    Operation_IFC mod_4308_inner <- mkFlatten(2);
    Operation_IFC mod_4308 <- mkDebugOperation(mod_4308_inner, "mod_4308");
    Operation_IFC mod_4309_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4309 <- mkDebugOperation(mod_4309_inner, "mod_4309");
    Broadcast_IFC#(4) mod_4310_inner <- mkBroadcast(4);
    Operation_IFC mod_4310 <- mkDebugOperation(mod_4310_inner.op, "mod_4310");
    PMU_IFC mod_4311_bufferize <- mkPMU(2);
    Operation_IFC mod_4311_inner = mod_4311_bufferize.operation;
    Operation_IFC mod_4311 <- mkDebugOperation(mod_4311_inner, "mod_4311");
    Broadcast_IFC#(2) mod_4312_inner <- mkBroadcast(2);
    Operation_IFC mod_4312 <- mkDebugOperation(mod_4312_inner.op, "mod_4312");
    PMU_IFC mod_4313_bufferize <- mkPMU(1);
    Operation_IFC mod_4313_inner = mod_4313_bufferize.operation;
    Operation_IFC mod_4313 <- mkDebugOperation(mod_4313_inner, "mod_4313");
    Operation_IFC mod_4314_inner <- mkBinaryMap(1051, matmul_t_tile);
    Operation_IFC mod_4314 <- mkDebugOperation(mod_4314_inner, "mod_4314");
    Operation_IFC mod_4315_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4315 <- mkDebugOperation(mod_4315_inner, "mod_4315");
    Operation_IFC mod_4316_inner <- mkBinaryMap(1819, mul_tile);
    Operation_IFC mod_4316 <- mkDebugOperation(mod_4316_inner, "mod_4316");
    PMU_IFC mod_4317_bufferize <- mkPMU(1);
    Operation_IFC mod_4317_inner = mod_4317_bufferize.operation;
    Operation_IFC mod_4317 <- mkDebugOperation(mod_4317_inner, "mod_4317");
    Operation_IFC mod_4318_inner <- mkBinaryMap(2353, matmul_t_tile);
    Operation_IFC mod_4318 <- mkDebugOperation(mod_4318_inner, "mod_4318");
    Operation_IFC mod_4319_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4319 <- mkDebugOperation(mod_4319_inner, "mod_4319");
    Operation_IFC mod_4320_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4320 <- mkDebugOperation(mod_4320_inner, "mod_4320");
    Operation_IFC mod_4321_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4321 <- mkDebugOperation(mod_4321_inner, "mod_4321");
    Operation_IFC mod_4322_inner <- mkBinaryMap(2718, mul_tile);
    Operation_IFC mod_4322 <- mkDebugOperation(mod_4322_inner, "mod_4322");
    PMU_IFC mod_4323_bufferize <- mkPMU(1);
    Operation_IFC mod_4323_inner = mod_4323_bufferize.operation;
    Operation_IFC mod_4323 <- mkDebugOperation(mod_4323_inner, "mod_4323");
    PMU_IFC mod_4324_bufferize <- mkPMU(2);
    Operation_IFC mod_4324_inner = mod_4324_bufferize.operation;
    Operation_IFC mod_4324 <- mkDebugOperation(mod_4324_inner, "mod_4324");
    PMU_IFC mod_4325_bufferize <- mkPMU(2);
    Operation_IFC mod_4325_inner = mod_4325_bufferize.operation;
    Operation_IFC mod_4325 <- mkDebugOperation(mod_4325_inner, "mod_4325");
    Operation_IFC mod_4326_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4326 <- mkDebugOperation(mod_4326_inner, "mod_4326");
    Operation_IFC mod_4327_inner <- mkFlatten(1);
    Operation_IFC mod_4327 <- mkDebugOperation(mod_4327_inner, "mod_4327");
    Operation_IFC mod_4328_inner <- mkFlatten(0);
    Operation_IFC mod_4328 <- mkDebugOperation(mod_4328_inner, "mod_4328");
    Operation_IFC mod_4329_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4329 <- mkDebugOperation(mod_4329_inner, "mod_4329");
    Operation_IFC mod_4330_inner <- mkUnaryMap(1691, silu_tile);
    Operation_IFC mod_4330 <- mkDebugOperation(mod_4330_inner, "mod_4330");
    Operation_IFC mod_4331_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4331 <- mkDebugOperation(mod_4331_inner, "mod_4331");
    Operation_IFC mod_4332_inner <- mkBinaryMap(1563, matmul_t_tile);
    Operation_IFC mod_4332 <- mkDebugOperation(mod_4332_inner, "mod_4332");
    PMU_IFC mod_4333_bufferize <- mkPMU(2);
    Operation_IFC mod_4333_inner = mod_4333_bufferize.operation;
    Operation_IFC mod_4333 <- mkDebugOperation(mod_4333_inner, "mod_4333");
    Operation_IFC mod_4334_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4334 <- mkDebugOperation(mod_4334_inner, "mod_4334");
    Operation_IFC mod_4335_inner <- mkFlatten(1);
    Operation_IFC mod_4335 <- mkDebugOperation(mod_4335_inner, "mod_4335");
    Operation_IFC mod_4336_inner <- mkFlatten(0);
    Operation_IFC mod_4336 <- mkDebugOperation(mod_4336_inner, "mod_4336");
    PMU_IFC mod_4337_bufferize <- mkPMU(1);
    Operation_IFC mod_4337_inner = mod_4337_bufferize.operation;
    Operation_IFC mod_4337 <- mkDebugOperation(mod_4337_inner, "mod_4337");
    Operation_IFC mod_4338_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4338 <- mkDebugOperation(mod_4338_inner, "mod_4338");
    PMU_IFC mod_4339_bufferize <- mkPMU(2);
    Operation_IFC mod_4339_inner = mod_4339_bufferize.operation;
    Operation_IFC mod_4339 <- mkDebugOperation(mod_4339_inner, "mod_4339");
    Operation_IFC mod_4340_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4340 <- mkDebugOperation(mod_4340_inner, "mod_4340");
    Operation_IFC mod_4341_inner <- mkFlatten(1);
    Operation_IFC mod_4341 <- mkDebugOperation(mod_4341_inner, "mod_4341");
    Operation_IFC mod_4342_inner <- mkFlatten(0);
    Operation_IFC mod_4342 <- mkDebugOperation(mod_4342_inner, "mod_4342");
    Operation_IFC mod_4343_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4343 <- mkDebugOperation(mod_4343_inner, "mod_4343");
    Operation_IFC mod_4344_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4344 <- mkDebugOperation(mod_4344_inner, "mod_4344");
    PMU_IFC mod_4345_bufferize <- mkPMU(2);
    Operation_IFC mod_4345_inner = mod_4345_bufferize.operation;
    Operation_IFC mod_4345 <- mkDebugOperation(mod_4345_inner, "mod_4345");
    rule rule_5566;
        ChannelMessage t;
        t <- mod_4343.get(0);
        mod_4313.put(1, t);
    endrule
    rule rule_5567;
        ChannelMessage t;
        t <- mod_4325.get(1);
        mod_4318.put(1, t);
    endrule
    rule rule_5568;
        ChannelMessage t;
        t <- mod_4313.get(0);
        mod_4343.put(0, t);
    endrule
    rule rule_5569;
        ChannelMessage t;
        t <- mod_4323.get(1);
        mod_4321.put(1, t);
    endrule
    rule rule_5570;
        ChannelMessage t;
        t <- mod_4332.get(0);
        mod_4331.put(0, t);
    endrule
    rule rule_5571;
        ChannelMessage t;
        t <- mod_4317.get(1);
        mod_4318.put(0, t);
    endrule
    rule rule_5572;
        ChannelMessage t;
        t <- mod_4321.get(1);
        mod_4322.put(1, t);
    endrule
    rule rule_5573;
        ChannelMessage t;
        t <- mod_4324.get(0);
        mod_4324.put(1, t);
    endrule
    rule rule_5574;
        ChannelMessage t;
        t <- mod_4316.get(0);
        mod_4317.put(0, t);
    endrule
    rule rule_5575;
        ChannelMessage t;
        t <- mod_4333.get(0);
        mod_4334.put(0, t);
    endrule
    rule rule_5576;
        ChannelMessage t;
        t <- mod_4341.get(0);
        mod_4339.put(0, t);
    endrule
    rule rule_5577;
        ChannelMessage t;
        t <- mod_4325.get(0);
        mod_4326.put(0, t);
    endrule
    rule rule_5578;
        ChannelMessage t;
        t <- mod_4328.get(0);
        mod_4327.put(0, t);
    endrule
    rule rule_5579;
        ChannelMessage t;
        t <- mod_4319.get(0);
        mod_4320.put(0, t);
    endrule
    rule rule_5580;
        ChannelMessage t;
        t <- mod_4333.get(1);
        mod_4332.put(1, t);
    endrule
    rule rule_5581;
        ChannelMessage t;
        t <- mod_4309.get(0);
        mod_4345.put(0, t);
    endrule
    rule rule_5582;
        ChannelMessage t;
        t <- mod_4334.get(0);
        mod_4333.put(1, t);
    endrule
    rule rule_5583;
        ChannelMessage t;
        t <- mod_4324.get(1);
        mod_4320.put(1, t);
    endrule
    rule rule_5584;
        ChannelMessage t;
        t <- mod_4327.get(0);
        mod_4325.put(0, t);
    endrule
    rule rule_5585;
        ChannelMessage t;
        t <- mod_4336.get(0);
        mod_4335.put(0, t);
    endrule
    rule rule_5586;
        ChannelMessage t;
        t <- mod_4337.get(0);
        mod_4338.put(0, t);
    endrule
    rule rule_5587;
        ChannelMessage t;
        t <- mod_4323.get(0);
        mod_4323.put(1, t);
    endrule
    rule rule_5588;
        ChannelMessage t;
        t <- mod_4311.get(1);
        mod_4312.put(0, t);
    endrule
    rule rule_5589;
        ChannelMessage t;
        t <- mod_4340.get(0);
        mod_4339.put(1, t);
    endrule
    rule rule_5590;
        ChannelMessage t;
        t <- mod_4337.get(1);
        mod_4332.put(0, t);
    endrule
    rule rule_5591;
        ChannelMessage t;
        t <- mod_4313.get(1);
        mod_4314.put(0, t);
    endrule
    rule rule_5592;
        ChannelMessage t;
        t <- mod_4345.get(1);
        mod_4309.put(1, t);
    endrule
    rule rule_5593;
        ChannelMessage t;
        t <- mod_4306.get(0);
        mod_4307.put(0, t);
    endrule
    rule rule_5594;
        ChannelMessage t;
        t <- mod_4335.get(0);
        mod_4333.put(0, t);
    endrule
    rule rule_5595;
        ChannelMessage t;
        t <- mod_4339.get(0);
        mod_4340.put(0, t);
    endrule
    rule rule_5596;
        ChannelMessage t;
        t <- mod_4311.get(0);
        mod_4344.put(0, t);
    endrule
    rule rule_5597;
        ChannelMessage t;
        t <- mod_4321.get(0);
        mod_4323.put(0, t);
    endrule
    rule rule_5598;
        ChannelMessage t;
        t <- mod_4326.get(0);
        mod_4325.put(1, t);
    endrule
    rule rule_5599;
        ChannelMessage t;
        t <- mod_4314.get(0);
        mod_4315.put(0, t);
    endrule
    rule rule_5600;
        ChannelMessage t;
        t <- mod_4342.get(0);
        mod_4341.put(0, t);
    endrule
    rule rule_5601;
        ChannelMessage t;
        t <- mod_4320.get(0);
        mod_4324.put(0, t);
    endrule
    rule rule_5602;
        ChannelMessage t;
        t <- mod_4320.get(1);
        mod_4321.put(0, t);
    endrule
    rule rule_5603;
        ChannelMessage t;
        t <- mod_4310.get(3);
        mod_4311.put(0, t);
    endrule
    rule rule_5604;
        ChannelMessage t;
        t <- mod_4312.get(1);
        mod_4313.put(0, t);
    endrule
    rule rule_5605;
        ChannelMessage t;
        t <- mod_4315.get(0);
        mod_4316.put(0, t);
    endrule
    rule rule_5606;
        ChannelMessage t;
        t <- mod_4309.get(1);
        mod_4310.put(0, t);
    endrule
    rule rule_5607;
        ChannelMessage t;
        t <- mod_4318.get(0);
        mod_4319.put(0, t);
    endrule
    rule rule_5608;
        ChannelMessage t;
        t <- mod_4308.get(0);
        mod_4309.put(0, t);
    endrule
    rule rule_5609;
        ChannelMessage t;
        t <- mod_4312.get(0);
        mod_4337.put(0, t);
    endrule
    rule rule_5610;
        ChannelMessage t;
        t <- mod_4329.get(0);
        mod_4317.put(1, t);
    endrule
    rule rule_5611;
        ChannelMessage t;
        t <- mod_4330.get(0);
        mod_4316.put(1, t);
    endrule
    rule rule_5612;
        ChannelMessage t;
        t <- mod_4331.get(0);
        mod_4330.put(0, t);
    endrule
    rule rule_5613;
        ChannelMessage t;
        t <- mod_4344.get(0);
        mod_4311.put(1, t);
    endrule
    rule rule_5614;
        ChannelMessage t;
        t <- mod_4338.get(0);
        mod_4337.put(1, t);
    endrule
    rule rule_5615;
        ChannelMessage t;
        t <- mod_4345.get(0);
        mod_4345.put(1, t);
    endrule
    rule rule_5616;
        ChannelMessage t;
        t <- mod_4307.get(0);
        mod_4308.put(0, t);
    endrule
    rule rule_5617;
        ChannelMessage t;
        t <- mod_4317.get(0);
        mod_4329.put(0, t);
    endrule
    rule rule_5618;
        ChannelMessage t;
        t <- mod_4339.get(1);
        mod_4314.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4306.put(0, t);
        end
        if (i == 1) begin
            mod_4322.put(0, t);
        end
        if (i == 2) begin
            mod_4328.put(0, t);
        end
        if (i == 3) begin
            mod_4336.put(0, t);
        end
        if (i == 4) begin
            mod_4342.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_4310.get(0);
        end
        if (i == 3) begin
            t <- mod_4310.get(1);
        end
        if (i == 2) begin
            t <- mod_4310.get(2);
        end
        if (i == 0) begin
            t <- mod_4322.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6140 (Operation_IFC);
    Operation_IFC mod_4347_inner <- mkReshape(2, 64);
    Operation_IFC mod_4347 <- mkDebugOperation(mod_4347_inner, "mod_4347");
    Operation_IFC mod_4348_inner <- mkFlatten(1);
    Operation_IFC mod_4348 <- mkDebugOperation(mod_4348_inner, "mod_4348");
    Operation_IFC mod_4349_inner <- mkFlatten(2);
    Operation_IFC mod_4349 <- mkDebugOperation(mod_4349_inner, "mod_4349");
    Operation_IFC mod_4350_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4350 <- mkDebugOperation(mod_4350_inner, "mod_4350");
    Broadcast_IFC#(4) mod_4351_inner <- mkBroadcast(4);
    Operation_IFC mod_4351 <- mkDebugOperation(mod_4351_inner.op, "mod_4351");
    PMU_IFC mod_4352_bufferize <- mkPMU(2);
    Operation_IFC mod_4352_inner = mod_4352_bufferize.operation;
    Operation_IFC mod_4352 <- mkDebugOperation(mod_4352_inner, "mod_4352");
    Broadcast_IFC#(2) mod_4353_inner <- mkBroadcast(2);
    Operation_IFC mod_4353 <- mkDebugOperation(mod_4353_inner.op, "mod_4353");
    PMU_IFC mod_4354_bufferize <- mkPMU(1);
    Operation_IFC mod_4354_inner = mod_4354_bufferize.operation;
    Operation_IFC mod_4354 <- mkDebugOperation(mod_4354_inner, "mod_4354");
    Operation_IFC mod_4355_inner <- mkBinaryMap(1050, matmul_t_tile);
    Operation_IFC mod_4355 <- mkDebugOperation(mod_4355_inner, "mod_4355");
    Operation_IFC mod_4356_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4356 <- mkDebugOperation(mod_4356_inner, "mod_4356");
    Operation_IFC mod_4357_inner <- mkBinaryMap(1818, mul_tile);
    Operation_IFC mod_4357 <- mkDebugOperation(mod_4357_inner, "mod_4357");
    PMU_IFC mod_4358_bufferize <- mkPMU(1);
    Operation_IFC mod_4358_inner = mod_4358_bufferize.operation;
    Operation_IFC mod_4358 <- mkDebugOperation(mod_4358_inner, "mod_4358");
    Operation_IFC mod_4359_inner <- mkBinaryMap(2351, matmul_t_tile);
    Operation_IFC mod_4359 <- mkDebugOperation(mod_4359_inner, "mod_4359");
    Operation_IFC mod_4360_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4360 <- mkDebugOperation(mod_4360_inner, "mod_4360");
    Operation_IFC mod_4361_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4361 <- mkDebugOperation(mod_4361_inner, "mod_4361");
    Operation_IFC mod_4362_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4362 <- mkDebugOperation(mod_4362_inner, "mod_4362");
    Operation_IFC mod_4363_inner <- mkBinaryMap(2717, mul_tile);
    Operation_IFC mod_4363 <- mkDebugOperation(mod_4363_inner, "mod_4363");
    PMU_IFC mod_4364_bufferize <- mkPMU(1);
    Operation_IFC mod_4364_inner = mod_4364_bufferize.operation;
    Operation_IFC mod_4364 <- mkDebugOperation(mod_4364_inner, "mod_4364");
    PMU_IFC mod_4365_bufferize <- mkPMU(2);
    Operation_IFC mod_4365_inner = mod_4365_bufferize.operation;
    Operation_IFC mod_4365 <- mkDebugOperation(mod_4365_inner, "mod_4365");
    PMU_IFC mod_4366_bufferize <- mkPMU(2);
    Operation_IFC mod_4366_inner = mod_4366_bufferize.operation;
    Operation_IFC mod_4366 <- mkDebugOperation(mod_4366_inner, "mod_4366");
    Operation_IFC mod_4367_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4367 <- mkDebugOperation(mod_4367_inner, "mod_4367");
    Operation_IFC mod_4368_inner <- mkFlatten(1);
    Operation_IFC mod_4368 <- mkDebugOperation(mod_4368_inner, "mod_4368");
    Operation_IFC mod_4369_inner <- mkFlatten(0);
    Operation_IFC mod_4369 <- mkDebugOperation(mod_4369_inner, "mod_4369");
    Operation_IFC mod_4370_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4370 <- mkDebugOperation(mod_4370_inner, "mod_4370");
    Operation_IFC mod_4371_inner <- mkUnaryMap(1690, silu_tile);
    Operation_IFC mod_4371 <- mkDebugOperation(mod_4371_inner, "mod_4371");
    Operation_IFC mod_4372_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4372 <- mkDebugOperation(mod_4372_inner, "mod_4372");
    Operation_IFC mod_4373_inner <- mkBinaryMap(1562, matmul_t_tile);
    Operation_IFC mod_4373 <- mkDebugOperation(mod_4373_inner, "mod_4373");
    PMU_IFC mod_4374_bufferize <- mkPMU(2);
    Operation_IFC mod_4374_inner = mod_4374_bufferize.operation;
    Operation_IFC mod_4374 <- mkDebugOperation(mod_4374_inner, "mod_4374");
    Operation_IFC mod_4375_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4375 <- mkDebugOperation(mod_4375_inner, "mod_4375");
    Operation_IFC mod_4376_inner <- mkFlatten(1);
    Operation_IFC mod_4376 <- mkDebugOperation(mod_4376_inner, "mod_4376");
    Operation_IFC mod_4377_inner <- mkFlatten(0);
    Operation_IFC mod_4377 <- mkDebugOperation(mod_4377_inner, "mod_4377");
    PMU_IFC mod_4378_bufferize <- mkPMU(1);
    Operation_IFC mod_4378_inner = mod_4378_bufferize.operation;
    Operation_IFC mod_4378 <- mkDebugOperation(mod_4378_inner, "mod_4378");
    Operation_IFC mod_4379_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4379 <- mkDebugOperation(mod_4379_inner, "mod_4379");
    PMU_IFC mod_4380_bufferize <- mkPMU(2);
    Operation_IFC mod_4380_inner = mod_4380_bufferize.operation;
    Operation_IFC mod_4380 <- mkDebugOperation(mod_4380_inner, "mod_4380");
    Operation_IFC mod_4381_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4381 <- mkDebugOperation(mod_4381_inner, "mod_4381");
    Operation_IFC mod_4382_inner <- mkFlatten(1);
    Operation_IFC mod_4382 <- mkDebugOperation(mod_4382_inner, "mod_4382");
    Operation_IFC mod_4383_inner <- mkFlatten(0);
    Operation_IFC mod_4383 <- mkDebugOperation(mod_4383_inner, "mod_4383");
    Operation_IFC mod_4384_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4384 <- mkDebugOperation(mod_4384_inner, "mod_4384");
    Operation_IFC mod_4385_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4385 <- mkDebugOperation(mod_4385_inner, "mod_4385");
    PMU_IFC mod_4386_bufferize <- mkPMU(2);
    Operation_IFC mod_4386_inner = mod_4386_bufferize.operation;
    Operation_IFC mod_4386 <- mkDebugOperation(mod_4386_inner, "mod_4386");
    rule rule_5619;
        ChannelMessage t;
        t <- mod_4350.get(0);
        mod_4386.put(0, t);
    endrule
    rule rule_5620;
        ChannelMessage t;
        t <- mod_4352.get(1);
        mod_4353.put(0, t);
    endrule
    rule rule_5621;
        ChannelMessage t;
        t <- mod_4383.get(0);
        mod_4382.put(0, t);
    endrule
    rule rule_5622;
        ChannelMessage t;
        t <- mod_4365.get(1);
        mod_4361.put(1, t);
    endrule
    rule rule_5623;
        ChannelMessage t;
        t <- mod_4361.get(1);
        mod_4362.put(0, t);
    endrule
    rule rule_5624;
        ChannelMessage t;
        t <- mod_4382.get(0);
        mod_4380.put(0, t);
    endrule
    rule rule_5625;
        ChannelMessage t;
        t <- mod_4348.get(0);
        mod_4349.put(0, t);
    endrule
    rule rule_5626;
        ChannelMessage t;
        t <- mod_4381.get(0);
        mod_4380.put(1, t);
    endrule
    rule rule_5627;
        ChannelMessage t;
        t <- mod_4385.get(0);
        mod_4352.put(1, t);
    endrule
    rule rule_5628;
        ChannelMessage t;
        t <- mod_4351.get(3);
        mod_4352.put(0, t);
    endrule
    rule rule_5629;
        ChannelMessage t;
        t <- mod_4386.get(0);
        mod_4386.put(1, t);
    endrule
    rule rule_5630;
        ChannelMessage t;
        t <- mod_4369.get(0);
        mod_4368.put(0, t);
    endrule
    rule rule_5631;
        ChannelMessage t;
        t <- mod_4355.get(0);
        mod_4356.put(0, t);
    endrule
    rule rule_5632;
        ChannelMessage t;
        t <- mod_4370.get(0);
        mod_4358.put(1, t);
    endrule
    rule rule_5633;
        ChannelMessage t;
        t <- mod_4364.get(1);
        mod_4362.put(1, t);
    endrule
    rule rule_5634;
        ChannelMessage t;
        t <- mod_4380.get(1);
        mod_4355.put(1, t);
    endrule
    rule rule_5635;
        ChannelMessage t;
        t <- mod_4384.get(0);
        mod_4354.put(1, t);
    endrule
    rule rule_5636;
        ChannelMessage t;
        t <- mod_4362.get(1);
        mod_4363.put(1, t);
    endrule
    rule rule_5637;
        ChannelMessage t;
        t <- mod_4372.get(0);
        mod_4371.put(0, t);
    endrule
    rule rule_5638;
        ChannelMessage t;
        t <- mod_4354.get(1);
        mod_4355.put(0, t);
    endrule
    rule rule_5639;
        ChannelMessage t;
        t <- mod_4353.get(1);
        mod_4354.put(0, t);
    endrule
    rule rule_5640;
        ChannelMessage t;
        t <- mod_4357.get(0);
        mod_4358.put(0, t);
    endrule
    rule rule_5641;
        ChannelMessage t;
        t <- mod_4358.get(1);
        mod_4359.put(0, t);
    endrule
    rule rule_5642;
        ChannelMessage t;
        t <- mod_4377.get(0);
        mod_4376.put(0, t);
    endrule
    rule rule_5643;
        ChannelMessage t;
        t <- mod_4366.get(0);
        mod_4367.put(0, t);
    endrule
    rule rule_5644;
        ChannelMessage t;
        t <- mod_4354.get(0);
        mod_4384.put(0, t);
    endrule
    rule rule_5645;
        ChannelMessage t;
        t <- mod_4350.get(1);
        mod_4351.put(0, t);
    endrule
    rule rule_5646;
        ChannelMessage t;
        t <- mod_4361.get(0);
        mod_4365.put(0, t);
    endrule
    rule rule_5647;
        ChannelMessage t;
        t <- mod_4358.get(0);
        mod_4370.put(0, t);
    endrule
    rule rule_5648;
        ChannelMessage t;
        t <- mod_4378.get(0);
        mod_4379.put(0, t);
    endrule
    rule rule_5649;
        ChannelMessage t;
        t <- mod_4365.get(0);
        mod_4365.put(1, t);
    endrule
    rule rule_5650;
        ChannelMessage t;
        t <- mod_4367.get(0);
        mod_4366.put(1, t);
    endrule
    rule rule_5651;
        ChannelMessage t;
        t <- mod_4368.get(0);
        mod_4366.put(0, t);
    endrule
    rule rule_5652;
        ChannelMessage t;
        t <- mod_4366.get(1);
        mod_4359.put(1, t);
    endrule
    rule rule_5653;
        ChannelMessage t;
        t <- mod_4373.get(0);
        mod_4372.put(0, t);
    endrule
    rule rule_5654;
        ChannelMessage t;
        t <- mod_4379.get(0);
        mod_4378.put(1, t);
    endrule
    rule rule_5655;
        ChannelMessage t;
        t <- mod_4380.get(0);
        mod_4381.put(0, t);
    endrule
    rule rule_5656;
        ChannelMessage t;
        t <- mod_4386.get(1);
        mod_4350.put(1, t);
    endrule
    rule rule_5657;
        ChannelMessage t;
        t <- mod_4378.get(1);
        mod_4373.put(0, t);
    endrule
    rule rule_5658;
        ChannelMessage t;
        t <- mod_4362.get(0);
        mod_4364.put(0, t);
    endrule
    rule rule_5659;
        ChannelMessage t;
        t <- mod_4374.get(0);
        mod_4375.put(0, t);
    endrule
    rule rule_5660;
        ChannelMessage t;
        t <- mod_4360.get(0);
        mod_4361.put(0, t);
    endrule
    rule rule_5661;
        ChannelMessage t;
        t <- mod_4374.get(1);
        mod_4373.put(1, t);
    endrule
    rule rule_5662;
        ChannelMessage t;
        t <- mod_4375.get(0);
        mod_4374.put(1, t);
    endrule
    rule rule_5663;
        ChannelMessage t;
        t <- mod_4364.get(0);
        mod_4364.put(1, t);
    endrule
    rule rule_5664;
        ChannelMessage t;
        t <- mod_4356.get(0);
        mod_4357.put(0, t);
    endrule
    rule rule_5665;
        ChannelMessage t;
        t <- mod_4371.get(0);
        mod_4357.put(1, t);
    endrule
    rule rule_5666;
        ChannelMessage t;
        t <- mod_4376.get(0);
        mod_4374.put(0, t);
    endrule
    rule rule_5667;
        ChannelMessage t;
        t <- mod_4353.get(0);
        mod_4378.put(0, t);
    endrule
    rule rule_5668;
        ChannelMessage t;
        t <- mod_4347.get(0);
        mod_4348.put(0, t);
    endrule
    rule rule_5669;
        ChannelMessage t;
        t <- mod_4349.get(0);
        mod_4350.put(0, t);
    endrule
    rule rule_5670;
        ChannelMessage t;
        t <- mod_4352.get(0);
        mod_4385.put(0, t);
    endrule
    rule rule_5671;
        ChannelMessage t;
        t <- mod_4359.get(0);
        mod_4360.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4347.put(0, t);
        end
        if (i == 1) begin
            mod_4363.put(0, t);
        end
        if (i == 2) begin
            mod_4369.put(0, t);
        end
        if (i == 3) begin
            mod_4377.put(0, t);
        end
        if (i == 4) begin
            mod_4383.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_4351.get(0);
        end
        if (i == 2) begin
            t <- mod_4351.get(1);
        end
        if (i == 3) begin
            t <- mod_4351.get(2);
        end
        if (i == 0) begin
            t <- mod_4363.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6141 (Operation_IFC);
    Operation_IFC mod_4388_inner <- mkReshape(2, 64);
    Operation_IFC mod_4388 <- mkDebugOperation(mod_4388_inner, "mod_4388");
    Operation_IFC mod_4389_inner <- mkFlatten(1);
    Operation_IFC mod_4389 <- mkDebugOperation(mod_4389_inner, "mod_4389");
    Operation_IFC mod_4390_inner <- mkFlatten(2);
    Operation_IFC mod_4390 <- mkDebugOperation(mod_4390_inner, "mod_4390");
    Operation_IFC mod_4391_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4391 <- mkDebugOperation(mod_4391_inner, "mod_4391");
    Broadcast_IFC#(4) mod_4392_inner <- mkBroadcast(4);
    Operation_IFC mod_4392 <- mkDebugOperation(mod_4392_inner.op, "mod_4392");
    PMU_IFC mod_4393_bufferize <- mkPMU(2);
    Operation_IFC mod_4393_inner = mod_4393_bufferize.operation;
    Operation_IFC mod_4393 <- mkDebugOperation(mod_4393_inner, "mod_4393");
    Broadcast_IFC#(2) mod_4394_inner <- mkBroadcast(2);
    Operation_IFC mod_4394 <- mkDebugOperation(mod_4394_inner.op, "mod_4394");
    PMU_IFC mod_4395_bufferize <- mkPMU(1);
    Operation_IFC mod_4395_inner = mod_4395_bufferize.operation;
    Operation_IFC mod_4395 <- mkDebugOperation(mod_4395_inner, "mod_4395");
    Operation_IFC mod_4396_inner <- mkBinaryMap(1049, matmul_t_tile);
    Operation_IFC mod_4396 <- mkDebugOperation(mod_4396_inner, "mod_4396");
    Operation_IFC mod_4397_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4397 <- mkDebugOperation(mod_4397_inner, "mod_4397");
    Operation_IFC mod_4398_inner <- mkBinaryMap(1817, mul_tile);
    Operation_IFC mod_4398 <- mkDebugOperation(mod_4398_inner, "mod_4398");
    PMU_IFC mod_4399_bufferize <- mkPMU(1);
    Operation_IFC mod_4399_inner = mod_4399_bufferize.operation;
    Operation_IFC mod_4399 <- mkDebugOperation(mod_4399_inner, "mod_4399");
    Operation_IFC mod_4400_inner <- mkBinaryMap(2349, matmul_t_tile);
    Operation_IFC mod_4400 <- mkDebugOperation(mod_4400_inner, "mod_4400");
    Operation_IFC mod_4401_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4401 <- mkDebugOperation(mod_4401_inner, "mod_4401");
    Operation_IFC mod_4402_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4402 <- mkDebugOperation(mod_4402_inner, "mod_4402");
    Operation_IFC mod_4403_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4403 <- mkDebugOperation(mod_4403_inner, "mod_4403");
    Operation_IFC mod_4404_inner <- mkBinaryMap(2716, mul_tile);
    Operation_IFC mod_4404 <- mkDebugOperation(mod_4404_inner, "mod_4404");
    PMU_IFC mod_4405_bufferize <- mkPMU(1);
    Operation_IFC mod_4405_inner = mod_4405_bufferize.operation;
    Operation_IFC mod_4405 <- mkDebugOperation(mod_4405_inner, "mod_4405");
    PMU_IFC mod_4406_bufferize <- mkPMU(2);
    Operation_IFC mod_4406_inner = mod_4406_bufferize.operation;
    Operation_IFC mod_4406 <- mkDebugOperation(mod_4406_inner, "mod_4406");
    PMU_IFC mod_4407_bufferize <- mkPMU(2);
    Operation_IFC mod_4407_inner = mod_4407_bufferize.operation;
    Operation_IFC mod_4407 <- mkDebugOperation(mod_4407_inner, "mod_4407");
    Operation_IFC mod_4408_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4408 <- mkDebugOperation(mod_4408_inner, "mod_4408");
    Operation_IFC mod_4409_inner <- mkFlatten(1);
    Operation_IFC mod_4409 <- mkDebugOperation(mod_4409_inner, "mod_4409");
    Operation_IFC mod_4410_inner <- mkFlatten(0);
    Operation_IFC mod_4410 <- mkDebugOperation(mod_4410_inner, "mod_4410");
    Operation_IFC mod_4411_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4411 <- mkDebugOperation(mod_4411_inner, "mod_4411");
    Operation_IFC mod_4412_inner <- mkUnaryMap(1689, silu_tile);
    Operation_IFC mod_4412 <- mkDebugOperation(mod_4412_inner, "mod_4412");
    Operation_IFC mod_4413_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4413 <- mkDebugOperation(mod_4413_inner, "mod_4413");
    Operation_IFC mod_4414_inner <- mkBinaryMap(1561, matmul_t_tile);
    Operation_IFC mod_4414 <- mkDebugOperation(mod_4414_inner, "mod_4414");
    PMU_IFC mod_4415_bufferize <- mkPMU(2);
    Operation_IFC mod_4415_inner = mod_4415_bufferize.operation;
    Operation_IFC mod_4415 <- mkDebugOperation(mod_4415_inner, "mod_4415");
    Operation_IFC mod_4416_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4416 <- mkDebugOperation(mod_4416_inner, "mod_4416");
    Operation_IFC mod_4417_inner <- mkFlatten(1);
    Operation_IFC mod_4417 <- mkDebugOperation(mod_4417_inner, "mod_4417");
    Operation_IFC mod_4418_inner <- mkFlatten(0);
    Operation_IFC mod_4418 <- mkDebugOperation(mod_4418_inner, "mod_4418");
    PMU_IFC mod_4419_bufferize <- mkPMU(1);
    Operation_IFC mod_4419_inner = mod_4419_bufferize.operation;
    Operation_IFC mod_4419 <- mkDebugOperation(mod_4419_inner, "mod_4419");
    Operation_IFC mod_4420_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4420 <- mkDebugOperation(mod_4420_inner, "mod_4420");
    PMU_IFC mod_4421_bufferize <- mkPMU(2);
    Operation_IFC mod_4421_inner = mod_4421_bufferize.operation;
    Operation_IFC mod_4421 <- mkDebugOperation(mod_4421_inner, "mod_4421");
    Operation_IFC mod_4422_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4422 <- mkDebugOperation(mod_4422_inner, "mod_4422");
    Operation_IFC mod_4423_inner <- mkFlatten(1);
    Operation_IFC mod_4423 <- mkDebugOperation(mod_4423_inner, "mod_4423");
    Operation_IFC mod_4424_inner <- mkFlatten(0);
    Operation_IFC mod_4424 <- mkDebugOperation(mod_4424_inner, "mod_4424");
    Operation_IFC mod_4425_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4425 <- mkDebugOperation(mod_4425_inner, "mod_4425");
    Operation_IFC mod_4426_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4426 <- mkDebugOperation(mod_4426_inner, "mod_4426");
    PMU_IFC mod_4427_bufferize <- mkPMU(2);
    Operation_IFC mod_4427_inner = mod_4427_bufferize.operation;
    Operation_IFC mod_4427 <- mkDebugOperation(mod_4427_inner, "mod_4427");
    rule rule_5672;
        ChannelMessage t;
        t <- mod_4400.get(0);
        mod_4401.put(0, t);
    endrule
    rule rule_5673;
        ChannelMessage t;
        t <- mod_4408.get(0);
        mod_4407.put(1, t);
    endrule
    rule rule_5674;
        ChannelMessage t;
        t <- mod_4406.get(0);
        mod_4406.put(1, t);
    endrule
    rule rule_5675;
        ChannelMessage t;
        t <- mod_4410.get(0);
        mod_4409.put(0, t);
    endrule
    rule rule_5676;
        ChannelMessage t;
        t <- mod_4389.get(0);
        mod_4390.put(0, t);
    endrule
    rule rule_5677;
        ChannelMessage t;
        t <- mod_4409.get(0);
        mod_4407.put(0, t);
    endrule
    rule rule_5678;
        ChannelMessage t;
        t <- mod_4393.get(1);
        mod_4394.put(0, t);
    endrule
    rule rule_5679;
        ChannelMessage t;
        t <- mod_4402.get(0);
        mod_4406.put(0, t);
    endrule
    rule rule_5680;
        ChannelMessage t;
        t <- mod_4399.get(1);
        mod_4400.put(0, t);
    endrule
    rule rule_5681;
        ChannelMessage t;
        t <- mod_4405.get(0);
        mod_4405.put(1, t);
    endrule
    rule rule_5682;
        ChannelMessage t;
        t <- mod_4406.get(1);
        mod_4402.put(1, t);
    endrule
    rule rule_5683;
        ChannelMessage t;
        t <- mod_4414.get(0);
        mod_4413.put(0, t);
    endrule
    rule rule_5684;
        ChannelMessage t;
        t <- mod_4392.get(3);
        mod_4393.put(0, t);
    endrule
    rule rule_5685;
        ChannelMessage t;
        t <- mod_4421.get(1);
        mod_4396.put(1, t);
    endrule
    rule rule_5686;
        ChannelMessage t;
        t <- mod_4401.get(0);
        mod_4402.put(0, t);
    endrule
    rule rule_5687;
        ChannelMessage t;
        t <- mod_4391.get(1);
        mod_4392.put(0, t);
    endrule
    rule rule_5688;
        ChannelMessage t;
        t <- mod_4415.get(0);
        mod_4416.put(0, t);
    endrule
    rule rule_5689;
        ChannelMessage t;
        t <- mod_4390.get(0);
        mod_4391.put(0, t);
    endrule
    rule rule_5690;
        ChannelMessage t;
        t <- mod_4398.get(0);
        mod_4399.put(0, t);
    endrule
    rule rule_5691;
        ChannelMessage t;
        t <- mod_4419.get(1);
        mod_4414.put(0, t);
    endrule
    rule rule_5692;
        ChannelMessage t;
        t <- mod_4396.get(0);
        mod_4397.put(0, t);
    endrule
    rule rule_5693;
        ChannelMessage t;
        t <- mod_4420.get(0);
        mod_4419.put(1, t);
    endrule
    rule rule_5694;
        ChannelMessage t;
        t <- mod_4399.get(0);
        mod_4411.put(0, t);
    endrule
    rule rule_5695;
        ChannelMessage t;
        t <- mod_4395.get(1);
        mod_4396.put(0, t);
    endrule
    rule rule_5696;
        ChannelMessage t;
        t <- mod_4394.get(1);
        mod_4395.put(0, t);
    endrule
    rule rule_5697;
        ChannelMessage t;
        t <- mod_4416.get(0);
        mod_4415.put(1, t);
    endrule
    rule rule_5698;
        ChannelMessage t;
        t <- mod_4424.get(0);
        mod_4423.put(0, t);
    endrule
    rule rule_5699;
        ChannelMessage t;
        t <- mod_4397.get(0);
        mod_4398.put(0, t);
    endrule
    rule rule_5700;
        ChannelMessage t;
        t <- mod_4425.get(0);
        mod_4395.put(1, t);
    endrule
    rule rule_5701;
        ChannelMessage t;
        t <- mod_4421.get(0);
        mod_4422.put(0, t);
    endrule
    rule rule_5702;
        ChannelMessage t;
        t <- mod_4417.get(0);
        mod_4415.put(0, t);
    endrule
    rule rule_5703;
        ChannelMessage t;
        t <- mod_4412.get(0);
        mod_4398.put(1, t);
    endrule
    rule rule_5704;
        ChannelMessage t;
        t <- mod_4405.get(1);
        mod_4403.put(1, t);
    endrule
    rule rule_5705;
        ChannelMessage t;
        t <- mod_4403.get(0);
        mod_4405.put(0, t);
    endrule
    rule rule_5706;
        ChannelMessage t;
        t <- mod_4407.get(0);
        mod_4408.put(0, t);
    endrule
    rule rule_5707;
        ChannelMessage t;
        t <- mod_4423.get(0);
        mod_4421.put(0, t);
    endrule
    rule rule_5708;
        ChannelMessage t;
        t <- mod_4426.get(0);
        mod_4393.put(1, t);
    endrule
    rule rule_5709;
        ChannelMessage t;
        t <- mod_4403.get(1);
        mod_4404.put(1, t);
    endrule
    rule rule_5710;
        ChannelMessage t;
        t <- mod_4427.get(1);
        mod_4391.put(1, t);
    endrule
    rule rule_5711;
        ChannelMessage t;
        t <- mod_4402.get(1);
        mod_4403.put(0, t);
    endrule
    rule rule_5712;
        ChannelMessage t;
        t <- mod_4418.get(0);
        mod_4417.put(0, t);
    endrule
    rule rule_5713;
        ChannelMessage t;
        t <- mod_4391.get(0);
        mod_4427.put(0, t);
    endrule
    rule rule_5714;
        ChannelMessage t;
        t <- mod_4413.get(0);
        mod_4412.put(0, t);
    endrule
    rule rule_5715;
        ChannelMessage t;
        t <- mod_4393.get(0);
        mod_4426.put(0, t);
    endrule
    rule rule_5716;
        ChannelMessage t;
        t <- mod_4419.get(0);
        mod_4420.put(0, t);
    endrule
    rule rule_5717;
        ChannelMessage t;
        t <- mod_4422.get(0);
        mod_4421.put(1, t);
    endrule
    rule rule_5718;
        ChannelMessage t;
        t <- mod_4395.get(0);
        mod_4425.put(0, t);
    endrule
    rule rule_5719;
        ChannelMessage t;
        t <- mod_4407.get(1);
        mod_4400.put(1, t);
    endrule
    rule rule_5720;
        ChannelMessage t;
        t <- mod_4427.get(0);
        mod_4427.put(1, t);
    endrule
    rule rule_5721;
        ChannelMessage t;
        t <- mod_4411.get(0);
        mod_4399.put(1, t);
    endrule
    rule rule_5722;
        ChannelMessage t;
        t <- mod_4415.get(1);
        mod_4414.put(1, t);
    endrule
    rule rule_5723;
        ChannelMessage t;
        t <- mod_4388.get(0);
        mod_4389.put(0, t);
    endrule
    rule rule_5724;
        ChannelMessage t;
        t <- mod_4394.get(0);
        mod_4419.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4388.put(0, t);
        end
        if (i == 1) begin
            mod_4404.put(0, t);
        end
        if (i == 2) begin
            mod_4410.put(0, t);
        end
        if (i == 3) begin
            mod_4418.put(0, t);
        end
        if (i == 4) begin
            mod_4424.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_4392.get(0);
        end
        if (i == 1) begin
            t <- mod_4392.get(1);
        end
        if (i == 2) begin
            t <- mod_4392.get(2);
        end
        if (i == 3) begin
            t <- mod_4404.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6142 (Operation_IFC);
    Operation_IFC mod_4429_inner <- mkReshape(2, 64);
    Operation_IFC mod_4429 <- mkDebugOperation(mod_4429_inner, "mod_4429");
    Operation_IFC mod_4430_inner <- mkFlatten(1);
    Operation_IFC mod_4430 <- mkDebugOperation(mod_4430_inner, "mod_4430");
    Operation_IFC mod_4431_inner <- mkFlatten(2);
    Operation_IFC mod_4431 <- mkDebugOperation(mod_4431_inner, "mod_4431");
    Operation_IFC mod_4432_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4432 <- mkDebugOperation(mod_4432_inner, "mod_4432");
    Broadcast_IFC#(4) mod_4433_inner <- mkBroadcast(4);
    Operation_IFC mod_4433 <- mkDebugOperation(mod_4433_inner.op, "mod_4433");
    PMU_IFC mod_4434_bufferize <- mkPMU(2);
    Operation_IFC mod_4434_inner = mod_4434_bufferize.operation;
    Operation_IFC mod_4434 <- mkDebugOperation(mod_4434_inner, "mod_4434");
    Broadcast_IFC#(2) mod_4435_inner <- mkBroadcast(2);
    Operation_IFC mod_4435 <- mkDebugOperation(mod_4435_inner.op, "mod_4435");
    PMU_IFC mod_4436_bufferize <- mkPMU(1);
    Operation_IFC mod_4436_inner = mod_4436_bufferize.operation;
    Operation_IFC mod_4436 <- mkDebugOperation(mod_4436_inner, "mod_4436");
    Operation_IFC mod_4437_inner <- mkBinaryMap(1048, matmul_t_tile);
    Operation_IFC mod_4437 <- mkDebugOperation(mod_4437_inner, "mod_4437");
    Operation_IFC mod_4438_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4438 <- mkDebugOperation(mod_4438_inner, "mod_4438");
    Operation_IFC mod_4439_inner <- mkBinaryMap(1816, mul_tile);
    Operation_IFC mod_4439 <- mkDebugOperation(mod_4439_inner, "mod_4439");
    PMU_IFC mod_4440_bufferize <- mkPMU(1);
    Operation_IFC mod_4440_inner = mod_4440_bufferize.operation;
    Operation_IFC mod_4440 <- mkDebugOperation(mod_4440_inner, "mod_4440");
    Operation_IFC mod_4441_inner <- mkBinaryMap(2347, matmul_t_tile);
    Operation_IFC mod_4441 <- mkDebugOperation(mod_4441_inner, "mod_4441");
    Operation_IFC mod_4442_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4442 <- mkDebugOperation(mod_4442_inner, "mod_4442");
    Operation_IFC mod_4443_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4443 <- mkDebugOperation(mod_4443_inner, "mod_4443");
    Operation_IFC mod_4444_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4444 <- mkDebugOperation(mod_4444_inner, "mod_4444");
    Operation_IFC mod_4445_inner <- mkBinaryMap(2715, mul_tile);
    Operation_IFC mod_4445 <- mkDebugOperation(mod_4445_inner, "mod_4445");
    PMU_IFC mod_4446_bufferize <- mkPMU(1);
    Operation_IFC mod_4446_inner = mod_4446_bufferize.operation;
    Operation_IFC mod_4446 <- mkDebugOperation(mod_4446_inner, "mod_4446");
    PMU_IFC mod_4447_bufferize <- mkPMU(2);
    Operation_IFC mod_4447_inner = mod_4447_bufferize.operation;
    Operation_IFC mod_4447 <- mkDebugOperation(mod_4447_inner, "mod_4447");
    PMU_IFC mod_4448_bufferize <- mkPMU(2);
    Operation_IFC mod_4448_inner = mod_4448_bufferize.operation;
    Operation_IFC mod_4448 <- mkDebugOperation(mod_4448_inner, "mod_4448");
    Operation_IFC mod_4449_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4449 <- mkDebugOperation(mod_4449_inner, "mod_4449");
    Operation_IFC mod_4450_inner <- mkFlatten(1);
    Operation_IFC mod_4450 <- mkDebugOperation(mod_4450_inner, "mod_4450");
    Operation_IFC mod_4451_inner <- mkFlatten(0);
    Operation_IFC mod_4451 <- mkDebugOperation(mod_4451_inner, "mod_4451");
    Operation_IFC mod_4452_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4452 <- mkDebugOperation(mod_4452_inner, "mod_4452");
    Operation_IFC mod_4453_inner <- mkUnaryMap(1688, silu_tile);
    Operation_IFC mod_4453 <- mkDebugOperation(mod_4453_inner, "mod_4453");
    Operation_IFC mod_4454_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4454 <- mkDebugOperation(mod_4454_inner, "mod_4454");
    Operation_IFC mod_4455_inner <- mkBinaryMap(1560, matmul_t_tile);
    Operation_IFC mod_4455 <- mkDebugOperation(mod_4455_inner, "mod_4455");
    PMU_IFC mod_4456_bufferize <- mkPMU(2);
    Operation_IFC mod_4456_inner = mod_4456_bufferize.operation;
    Operation_IFC mod_4456 <- mkDebugOperation(mod_4456_inner, "mod_4456");
    Operation_IFC mod_4457_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4457 <- mkDebugOperation(mod_4457_inner, "mod_4457");
    Operation_IFC mod_4458_inner <- mkFlatten(1);
    Operation_IFC mod_4458 <- mkDebugOperation(mod_4458_inner, "mod_4458");
    Operation_IFC mod_4459_inner <- mkFlatten(0);
    Operation_IFC mod_4459 <- mkDebugOperation(mod_4459_inner, "mod_4459");
    PMU_IFC mod_4460_bufferize <- mkPMU(1);
    Operation_IFC mod_4460_inner = mod_4460_bufferize.operation;
    Operation_IFC mod_4460 <- mkDebugOperation(mod_4460_inner, "mod_4460");
    Operation_IFC mod_4461_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4461 <- mkDebugOperation(mod_4461_inner, "mod_4461");
    PMU_IFC mod_4462_bufferize <- mkPMU(2);
    Operation_IFC mod_4462_inner = mod_4462_bufferize.operation;
    Operation_IFC mod_4462 <- mkDebugOperation(mod_4462_inner, "mod_4462");
    Operation_IFC mod_4463_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4463 <- mkDebugOperation(mod_4463_inner, "mod_4463");
    Operation_IFC mod_4464_inner <- mkFlatten(1);
    Operation_IFC mod_4464 <- mkDebugOperation(mod_4464_inner, "mod_4464");
    Operation_IFC mod_4465_inner <- mkFlatten(0);
    Operation_IFC mod_4465 <- mkDebugOperation(mod_4465_inner, "mod_4465");
    Operation_IFC mod_4466_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4466 <- mkDebugOperation(mod_4466_inner, "mod_4466");
    Operation_IFC mod_4467_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4467 <- mkDebugOperation(mod_4467_inner, "mod_4467");
    PMU_IFC mod_4468_bufferize <- mkPMU(2);
    Operation_IFC mod_4468_inner = mod_4468_bufferize.operation;
    Operation_IFC mod_4468 <- mkDebugOperation(mod_4468_inner, "mod_4468");
    rule rule_5725;
        ChannelMessage t;
        t <- mod_4444.get(0);
        mod_4446.put(0, t);
    endrule
    rule rule_5726;
        ChannelMessage t;
        t <- mod_4455.get(0);
        mod_4454.put(0, t);
    endrule
    rule rule_5727;
        ChannelMessage t;
        t <- mod_4431.get(0);
        mod_4432.put(0, t);
    endrule
    rule rule_5728;
        ChannelMessage t;
        t <- mod_4433.get(3);
        mod_4434.put(0, t);
    endrule
    rule rule_5729;
        ChannelMessage t;
        t <- mod_4456.get(0);
        mod_4457.put(0, t);
    endrule
    rule rule_5730;
        ChannelMessage t;
        t <- mod_4458.get(0);
        mod_4456.put(0, t);
    endrule
    rule rule_5731;
        ChannelMessage t;
        t <- mod_4464.get(0);
        mod_4462.put(0, t);
    endrule
    rule rule_5732;
        ChannelMessage t;
        t <- mod_4446.get(0);
        mod_4446.put(1, t);
    endrule
    rule rule_5733;
        ChannelMessage t;
        t <- mod_4429.get(0);
        mod_4430.put(0, t);
    endrule
    rule rule_5734;
        ChannelMessage t;
        t <- mod_4448.get(0);
        mod_4449.put(0, t);
    endrule
    rule rule_5735;
        ChannelMessage t;
        t <- mod_4466.get(0);
        mod_4436.put(1, t);
    endrule
    rule rule_5736;
        ChannelMessage t;
        t <- mod_4434.get(0);
        mod_4467.put(0, t);
    endrule
    rule rule_5737;
        ChannelMessage t;
        t <- mod_4468.get(1);
        mod_4432.put(1, t);
    endrule
    rule rule_5738;
        ChannelMessage t;
        t <- mod_4452.get(0);
        mod_4440.put(1, t);
    endrule
    rule rule_5739;
        ChannelMessage t;
        t <- mod_4444.get(1);
        mod_4445.put(1, t);
    endrule
    rule rule_5740;
        ChannelMessage t;
        t <- mod_4459.get(0);
        mod_4458.put(0, t);
    endrule
    rule rule_5741;
        ChannelMessage t;
        t <- mod_4462.get(1);
        mod_4437.put(1, t);
    endrule
    rule rule_5742;
        ChannelMessage t;
        t <- mod_4443.get(0);
        mod_4447.put(0, t);
    endrule
    rule rule_5743;
        ChannelMessage t;
        t <- mod_4440.get(1);
        mod_4441.put(0, t);
    endrule
    rule rule_5744;
        ChannelMessage t;
        t <- mod_4461.get(0);
        mod_4460.put(1, t);
    endrule
    rule rule_5745;
        ChannelMessage t;
        t <- mod_4432.get(0);
        mod_4468.put(0, t);
    endrule
    rule rule_5746;
        ChannelMessage t;
        t <- mod_4446.get(1);
        mod_4444.put(1, t);
    endrule
    rule rule_5747;
        ChannelMessage t;
        t <- mod_4460.get(0);
        mod_4461.put(0, t);
    endrule
    rule rule_5748;
        ChannelMessage t;
        t <- mod_4449.get(0);
        mod_4448.put(1, t);
    endrule
    rule rule_5749;
        ChannelMessage t;
        t <- mod_4437.get(0);
        mod_4438.put(0, t);
    endrule
    rule rule_5750;
        ChannelMessage t;
        t <- mod_4462.get(0);
        mod_4463.put(0, t);
    endrule
    rule rule_5751;
        ChannelMessage t;
        t <- mod_4465.get(0);
        mod_4464.put(0, t);
    endrule
    rule rule_5752;
        ChannelMessage t;
        t <- mod_4453.get(0);
        mod_4439.put(1, t);
    endrule
    rule rule_5753;
        ChannelMessage t;
        t <- mod_4435.get(1);
        mod_4436.put(0, t);
    endrule
    rule rule_5754;
        ChannelMessage t;
        t <- mod_4438.get(0);
        mod_4439.put(0, t);
    endrule
    rule rule_5755;
        ChannelMessage t;
        t <- mod_4441.get(0);
        mod_4442.put(0, t);
    endrule
    rule rule_5756;
        ChannelMessage t;
        t <- mod_4457.get(0);
        mod_4456.put(1, t);
    endrule
    rule rule_5757;
        ChannelMessage t;
        t <- mod_4432.get(1);
        mod_4433.put(0, t);
    endrule
    rule rule_5758;
        ChannelMessage t;
        t <- mod_4450.get(0);
        mod_4448.put(0, t);
    endrule
    rule rule_5759;
        ChannelMessage t;
        t <- mod_4456.get(1);
        mod_4455.put(1, t);
    endrule
    rule rule_5760;
        ChannelMessage t;
        t <- mod_4436.get(0);
        mod_4466.put(0, t);
    endrule
    rule rule_5761;
        ChannelMessage t;
        t <- mod_4451.get(0);
        mod_4450.put(0, t);
    endrule
    rule rule_5762;
        ChannelMessage t;
        t <- mod_4443.get(1);
        mod_4444.put(0, t);
    endrule
    rule rule_5763;
        ChannelMessage t;
        t <- mod_4460.get(1);
        mod_4455.put(0, t);
    endrule
    rule rule_5764;
        ChannelMessage t;
        t <- mod_4447.get(1);
        mod_4443.put(1, t);
    endrule
    rule rule_5765;
        ChannelMessage t;
        t <- mod_4442.get(0);
        mod_4443.put(0, t);
    endrule
    rule rule_5766;
        ChannelMessage t;
        t <- mod_4440.get(0);
        mod_4452.put(0, t);
    endrule
    rule rule_5767;
        ChannelMessage t;
        t <- mod_4448.get(1);
        mod_4441.put(1, t);
    endrule
    rule rule_5768;
        ChannelMessage t;
        t <- mod_4454.get(0);
        mod_4453.put(0, t);
    endrule
    rule rule_5769;
        ChannelMessage t;
        t <- mod_4447.get(0);
        mod_4447.put(1, t);
    endrule
    rule rule_5770;
        ChannelMessage t;
        t <- mod_4468.get(0);
        mod_4468.put(1, t);
    endrule
    rule rule_5771;
        ChannelMessage t;
        t <- mod_4467.get(0);
        mod_4434.put(1, t);
    endrule
    rule rule_5772;
        ChannelMessage t;
        t <- mod_4439.get(0);
        mod_4440.put(0, t);
    endrule
    rule rule_5773;
        ChannelMessage t;
        t <- mod_4434.get(1);
        mod_4435.put(0, t);
    endrule
    rule rule_5774;
        ChannelMessage t;
        t <- mod_4436.get(1);
        mod_4437.put(0, t);
    endrule
    rule rule_5775;
        ChannelMessage t;
        t <- mod_4435.get(0);
        mod_4460.put(0, t);
    endrule
    rule rule_5776;
        ChannelMessage t;
        t <- mod_4430.get(0);
        mod_4431.put(0, t);
    endrule
    rule rule_5777;
        ChannelMessage t;
        t <- mod_4463.get(0);
        mod_4462.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4429.put(0, t);
        end
        if (i == 1) begin
            mod_4445.put(0, t);
        end
        if (i == 2) begin
            mod_4451.put(0, t);
        end
        if (i == 3) begin
            mod_4459.put(0, t);
        end
        if (i == 4) begin
            mod_4465.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_4433.get(0);
        end
        if (i == 1) begin
            t <- mod_4433.get(1);
        end
        if (i == 3) begin
            t <- mod_4433.get(2);
        end
        if (i == 2) begin
            t <- mod_4445.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6143 (Operation_IFC);
    Operation_IFC mod_4470_inner <- mkReshape(2, 64);
    Operation_IFC mod_4470 <- mkDebugOperation(mod_4470_inner, "mod_4470");
    Operation_IFC mod_4471_inner <- mkFlatten(1);
    Operation_IFC mod_4471 <- mkDebugOperation(mod_4471_inner, "mod_4471");
    Operation_IFC mod_4472_inner <- mkFlatten(2);
    Operation_IFC mod_4472 <- mkDebugOperation(mod_4472_inner, "mod_4472");
    Operation_IFC mod_4473_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4473 <- mkDebugOperation(mod_4473_inner, "mod_4473");
    Broadcast_IFC#(4) mod_4474_inner <- mkBroadcast(4);
    Operation_IFC mod_4474 <- mkDebugOperation(mod_4474_inner.op, "mod_4474");
    PMU_IFC mod_4475_bufferize <- mkPMU(2);
    Operation_IFC mod_4475_inner = mod_4475_bufferize.operation;
    Operation_IFC mod_4475 <- mkDebugOperation(mod_4475_inner, "mod_4475");
    Broadcast_IFC#(2) mod_4476_inner <- mkBroadcast(2);
    Operation_IFC mod_4476 <- mkDebugOperation(mod_4476_inner.op, "mod_4476");
    PMU_IFC mod_4477_bufferize <- mkPMU(1);
    Operation_IFC mod_4477_inner = mod_4477_bufferize.operation;
    Operation_IFC mod_4477 <- mkDebugOperation(mod_4477_inner, "mod_4477");
    Operation_IFC mod_4478_inner <- mkBinaryMap(1047, matmul_t_tile);
    Operation_IFC mod_4478 <- mkDebugOperation(mod_4478_inner, "mod_4478");
    Operation_IFC mod_4479_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4479 <- mkDebugOperation(mod_4479_inner, "mod_4479");
    Operation_IFC mod_4480_inner <- mkBinaryMap(1815, mul_tile);
    Operation_IFC mod_4480 <- mkDebugOperation(mod_4480_inner, "mod_4480");
    PMU_IFC mod_4481_bufferize <- mkPMU(1);
    Operation_IFC mod_4481_inner = mod_4481_bufferize.operation;
    Operation_IFC mod_4481 <- mkDebugOperation(mod_4481_inner, "mod_4481");
    Operation_IFC mod_4482_inner <- mkBinaryMap(2345, matmul_t_tile);
    Operation_IFC mod_4482 <- mkDebugOperation(mod_4482_inner, "mod_4482");
    Operation_IFC mod_4483_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4483 <- mkDebugOperation(mod_4483_inner, "mod_4483");
    Operation_IFC mod_4484_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4484 <- mkDebugOperation(mod_4484_inner, "mod_4484");
    Operation_IFC mod_4485_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4485 <- mkDebugOperation(mod_4485_inner, "mod_4485");
    Operation_IFC mod_4486_inner <- mkBinaryMap(2714, mul_tile);
    Operation_IFC mod_4486 <- mkDebugOperation(mod_4486_inner, "mod_4486");
    PMU_IFC mod_4487_bufferize <- mkPMU(1);
    Operation_IFC mod_4487_inner = mod_4487_bufferize.operation;
    Operation_IFC mod_4487 <- mkDebugOperation(mod_4487_inner, "mod_4487");
    PMU_IFC mod_4488_bufferize <- mkPMU(2);
    Operation_IFC mod_4488_inner = mod_4488_bufferize.operation;
    Operation_IFC mod_4488 <- mkDebugOperation(mod_4488_inner, "mod_4488");
    PMU_IFC mod_4489_bufferize <- mkPMU(2);
    Operation_IFC mod_4489_inner = mod_4489_bufferize.operation;
    Operation_IFC mod_4489 <- mkDebugOperation(mod_4489_inner, "mod_4489");
    Operation_IFC mod_4490_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4490 <- mkDebugOperation(mod_4490_inner, "mod_4490");
    Operation_IFC mod_4491_inner <- mkFlatten(1);
    Operation_IFC mod_4491 <- mkDebugOperation(mod_4491_inner, "mod_4491");
    Operation_IFC mod_4492_inner <- mkFlatten(0);
    Operation_IFC mod_4492 <- mkDebugOperation(mod_4492_inner, "mod_4492");
    Operation_IFC mod_4493_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4493 <- mkDebugOperation(mod_4493_inner, "mod_4493");
    Operation_IFC mod_4494_inner <- mkUnaryMap(1687, silu_tile);
    Operation_IFC mod_4494 <- mkDebugOperation(mod_4494_inner, "mod_4494");
    Operation_IFC mod_4495_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4495 <- mkDebugOperation(mod_4495_inner, "mod_4495");
    Operation_IFC mod_4496_inner <- mkBinaryMap(1559, matmul_t_tile);
    Operation_IFC mod_4496 <- mkDebugOperation(mod_4496_inner, "mod_4496");
    PMU_IFC mod_4497_bufferize <- mkPMU(2);
    Operation_IFC mod_4497_inner = mod_4497_bufferize.operation;
    Operation_IFC mod_4497 <- mkDebugOperation(mod_4497_inner, "mod_4497");
    Operation_IFC mod_4498_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4498 <- mkDebugOperation(mod_4498_inner, "mod_4498");
    Operation_IFC mod_4499_inner <- mkFlatten(1);
    Operation_IFC mod_4499 <- mkDebugOperation(mod_4499_inner, "mod_4499");
    Operation_IFC mod_4500_inner <- mkFlatten(0);
    Operation_IFC mod_4500 <- mkDebugOperation(mod_4500_inner, "mod_4500");
    PMU_IFC mod_4501_bufferize <- mkPMU(1);
    Operation_IFC mod_4501_inner = mod_4501_bufferize.operation;
    Operation_IFC mod_4501 <- mkDebugOperation(mod_4501_inner, "mod_4501");
    Operation_IFC mod_4502_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4502 <- mkDebugOperation(mod_4502_inner, "mod_4502");
    PMU_IFC mod_4503_bufferize <- mkPMU(2);
    Operation_IFC mod_4503_inner = mod_4503_bufferize.operation;
    Operation_IFC mod_4503 <- mkDebugOperation(mod_4503_inner, "mod_4503");
    Operation_IFC mod_4504_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4504 <- mkDebugOperation(mod_4504_inner, "mod_4504");
    Operation_IFC mod_4505_inner <- mkFlatten(1);
    Operation_IFC mod_4505 <- mkDebugOperation(mod_4505_inner, "mod_4505");
    Operation_IFC mod_4506_inner <- mkFlatten(0);
    Operation_IFC mod_4506 <- mkDebugOperation(mod_4506_inner, "mod_4506");
    Operation_IFC mod_4507_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4507 <- mkDebugOperation(mod_4507_inner, "mod_4507");
    Operation_IFC mod_4508_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4508 <- mkDebugOperation(mod_4508_inner, "mod_4508");
    PMU_IFC mod_4509_bufferize <- mkPMU(2);
    Operation_IFC mod_4509_inner = mod_4509_bufferize.operation;
    Operation_IFC mod_4509 <- mkDebugOperation(mod_4509_inner, "mod_4509");
    rule rule_5778;
        ChannelMessage t;
        t <- mod_4497.get(1);
        mod_4496.put(1, t);
    endrule
    rule rule_5779;
        ChannelMessage t;
        t <- mod_4501.get(0);
        mod_4502.put(0, t);
    endrule
    rule rule_5780;
        ChannelMessage t;
        t <- mod_4470.get(0);
        mod_4471.put(0, t);
    endrule
    rule rule_5781;
        ChannelMessage t;
        t <- mod_4503.get(0);
        mod_4504.put(0, t);
    endrule
    rule rule_5782;
        ChannelMessage t;
        t <- mod_4472.get(0);
        mod_4473.put(0, t);
    endrule
    rule rule_5783;
        ChannelMessage t;
        t <- mod_4477.get(0);
        mod_4507.put(0, t);
    endrule
    rule rule_5784;
        ChannelMessage t;
        t <- mod_4509.get(0);
        mod_4509.put(1, t);
    endrule
    rule rule_5785;
        ChannelMessage t;
        t <- mod_4501.get(1);
        mod_4496.put(0, t);
    endrule
    rule rule_5786;
        ChannelMessage t;
        t <- mod_4476.get(1);
        mod_4477.put(0, t);
    endrule
    rule rule_5787;
        ChannelMessage t;
        t <- mod_4492.get(0);
        mod_4491.put(0, t);
    endrule
    rule rule_5788;
        ChannelMessage t;
        t <- mod_4473.get(1);
        mod_4474.put(0, t);
    endrule
    rule rule_5789;
        ChannelMessage t;
        t <- mod_4475.get(1);
        mod_4476.put(0, t);
    endrule
    rule rule_5790;
        ChannelMessage t;
        t <- mod_4481.get(0);
        mod_4493.put(0, t);
    endrule
    rule rule_5791;
        ChannelMessage t;
        t <- mod_4481.get(1);
        mod_4482.put(0, t);
    endrule
    rule rule_5792;
        ChannelMessage t;
        t <- mod_4498.get(0);
        mod_4497.put(1, t);
    endrule
    rule rule_5793;
        ChannelMessage t;
        t <- mod_4508.get(0);
        mod_4475.put(1, t);
    endrule
    rule rule_5794;
        ChannelMessage t;
        t <- mod_4491.get(0);
        mod_4489.put(0, t);
    endrule
    rule rule_5795;
        ChannelMessage t;
        t <- mod_4489.get(1);
        mod_4482.put(1, t);
    endrule
    rule rule_5796;
        ChannelMessage t;
        t <- mod_4493.get(0);
        mod_4481.put(1, t);
    endrule
    rule rule_5797;
        ChannelMessage t;
        t <- mod_4504.get(0);
        mod_4503.put(1, t);
    endrule
    rule rule_5798;
        ChannelMessage t;
        t <- mod_4485.get(0);
        mod_4487.put(0, t);
    endrule
    rule rule_5799;
        ChannelMessage t;
        t <- mod_4507.get(0);
        mod_4477.put(1, t);
    endrule
    rule rule_5800;
        ChannelMessage t;
        t <- mod_4494.get(0);
        mod_4480.put(1, t);
    endrule
    rule rule_5801;
        ChannelMessage t;
        t <- mod_4480.get(0);
        mod_4481.put(0, t);
    endrule
    rule rule_5802;
        ChannelMessage t;
        t <- mod_4487.get(1);
        mod_4485.put(1, t);
    endrule
    rule rule_5803;
        ChannelMessage t;
        t <- mod_4482.get(0);
        mod_4483.put(0, t);
    endrule
    rule rule_5804;
        ChannelMessage t;
        t <- mod_4505.get(0);
        mod_4503.put(0, t);
    endrule
    rule rule_5805;
        ChannelMessage t;
        t <- mod_4474.get(3);
        mod_4475.put(0, t);
    endrule
    rule rule_5806;
        ChannelMessage t;
        t <- mod_4471.get(0);
        mod_4472.put(0, t);
    endrule
    rule rule_5807;
        ChannelMessage t;
        t <- mod_4485.get(1);
        mod_4486.put(1, t);
    endrule
    rule rule_5808;
        ChannelMessage t;
        t <- mod_4487.get(0);
        mod_4487.put(1, t);
    endrule
    rule rule_5809;
        ChannelMessage t;
        t <- mod_4502.get(0);
        mod_4501.put(1, t);
    endrule
    rule rule_5810;
        ChannelMessage t;
        t <- mod_4479.get(0);
        mod_4480.put(0, t);
    endrule
    rule rule_5811;
        ChannelMessage t;
        t <- mod_4499.get(0);
        mod_4497.put(0, t);
    endrule
    rule rule_5812;
        ChannelMessage t;
        t <- mod_4484.get(0);
        mod_4488.put(0, t);
    endrule
    rule rule_5813;
        ChannelMessage t;
        t <- mod_4483.get(0);
        mod_4484.put(0, t);
    endrule
    rule rule_5814;
        ChannelMessage t;
        t <- mod_4484.get(1);
        mod_4485.put(0, t);
    endrule
    rule rule_5815;
        ChannelMessage t;
        t <- mod_4490.get(0);
        mod_4489.put(1, t);
    endrule
    rule rule_5816;
        ChannelMessage t;
        t <- mod_4473.get(0);
        mod_4509.put(0, t);
    endrule
    rule rule_5817;
        ChannelMessage t;
        t <- mod_4495.get(0);
        mod_4494.put(0, t);
    endrule
    rule rule_5818;
        ChannelMessage t;
        t <- mod_4488.get(1);
        mod_4484.put(1, t);
    endrule
    rule rule_5819;
        ChannelMessage t;
        t <- mod_4506.get(0);
        mod_4505.put(0, t);
    endrule
    rule rule_5820;
        ChannelMessage t;
        t <- mod_4496.get(0);
        mod_4495.put(0, t);
    endrule
    rule rule_5821;
        ChannelMessage t;
        t <- mod_4476.get(0);
        mod_4501.put(0, t);
    endrule
    rule rule_5822;
        ChannelMessage t;
        t <- mod_4478.get(0);
        mod_4479.put(0, t);
    endrule
    rule rule_5823;
        ChannelMessage t;
        t <- mod_4488.get(0);
        mod_4488.put(1, t);
    endrule
    rule rule_5824;
        ChannelMessage t;
        t <- mod_4489.get(0);
        mod_4490.put(0, t);
    endrule
    rule rule_5825;
        ChannelMessage t;
        t <- mod_4500.get(0);
        mod_4499.put(0, t);
    endrule
    rule rule_5826;
        ChannelMessage t;
        t <- mod_4503.get(1);
        mod_4478.put(1, t);
    endrule
    rule rule_5827;
        ChannelMessage t;
        t <- mod_4475.get(0);
        mod_4508.put(0, t);
    endrule
    rule rule_5828;
        ChannelMessage t;
        t <- mod_4477.get(1);
        mod_4478.put(0, t);
    endrule
    rule rule_5829;
        ChannelMessage t;
        t <- mod_4497.get(0);
        mod_4498.put(0, t);
    endrule
    rule rule_5830;
        ChannelMessage t;
        t <- mod_4509.get(1);
        mod_4473.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4470.put(0, t);
        end
        if (i == 1) begin
            mod_4486.put(0, t);
        end
        if (i == 2) begin
            mod_4492.put(0, t);
        end
        if (i == 3) begin
            mod_4500.put(0, t);
        end
        if (i == 4) begin
            mod_4506.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_4474.get(0);
        end
        if (i == 2) begin
            t <- mod_4474.get(1);
        end
        if (i == 1) begin
            t <- mod_4474.get(2);
        end
        if (i == 3) begin
            t <- mod_4486.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6144 (Operation_IFC);
    Operation_IFC mod_4511_inner <- mkReshape(2, 64);
    Operation_IFC mod_4511 <- mkDebugOperation(mod_4511_inner, "mod_4511");
    Operation_IFC mod_4512_inner <- mkFlatten(1);
    Operation_IFC mod_4512 <- mkDebugOperation(mod_4512_inner, "mod_4512");
    Operation_IFC mod_4513_inner <- mkFlatten(2);
    Operation_IFC mod_4513 <- mkDebugOperation(mod_4513_inner, "mod_4513");
    Operation_IFC mod_4514_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4514 <- mkDebugOperation(mod_4514_inner, "mod_4514");
    Broadcast_IFC#(4) mod_4515_inner <- mkBroadcast(4);
    Operation_IFC mod_4515 <- mkDebugOperation(mod_4515_inner.op, "mod_4515");
    PMU_IFC mod_4516_bufferize <- mkPMU(2);
    Operation_IFC mod_4516_inner = mod_4516_bufferize.operation;
    Operation_IFC mod_4516 <- mkDebugOperation(mod_4516_inner, "mod_4516");
    Broadcast_IFC#(2) mod_4517_inner <- mkBroadcast(2);
    Operation_IFC mod_4517 <- mkDebugOperation(mod_4517_inner.op, "mod_4517");
    PMU_IFC mod_4518_bufferize <- mkPMU(1);
    Operation_IFC mod_4518_inner = mod_4518_bufferize.operation;
    Operation_IFC mod_4518 <- mkDebugOperation(mod_4518_inner, "mod_4518");
    Operation_IFC mod_4519_inner <- mkBinaryMap(1046, matmul_t_tile);
    Operation_IFC mod_4519 <- mkDebugOperation(mod_4519_inner, "mod_4519");
    Operation_IFC mod_4520_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4520 <- mkDebugOperation(mod_4520_inner, "mod_4520");
    Operation_IFC mod_4521_inner <- mkBinaryMap(1814, mul_tile);
    Operation_IFC mod_4521 <- mkDebugOperation(mod_4521_inner, "mod_4521");
    PMU_IFC mod_4522_bufferize <- mkPMU(1);
    Operation_IFC mod_4522_inner = mod_4522_bufferize.operation;
    Operation_IFC mod_4522 <- mkDebugOperation(mod_4522_inner, "mod_4522");
    Operation_IFC mod_4523_inner <- mkBinaryMap(2343, matmul_t_tile);
    Operation_IFC mod_4523 <- mkDebugOperation(mod_4523_inner, "mod_4523");
    Operation_IFC mod_4524_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4524 <- mkDebugOperation(mod_4524_inner, "mod_4524");
    Operation_IFC mod_4525_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4525 <- mkDebugOperation(mod_4525_inner, "mod_4525");
    Operation_IFC mod_4526_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4526 <- mkDebugOperation(mod_4526_inner, "mod_4526");
    Operation_IFC mod_4527_inner <- mkBinaryMap(2713, mul_tile);
    Operation_IFC mod_4527 <- mkDebugOperation(mod_4527_inner, "mod_4527");
    PMU_IFC mod_4528_bufferize <- mkPMU(1);
    Operation_IFC mod_4528_inner = mod_4528_bufferize.operation;
    Operation_IFC mod_4528 <- mkDebugOperation(mod_4528_inner, "mod_4528");
    PMU_IFC mod_4529_bufferize <- mkPMU(2);
    Operation_IFC mod_4529_inner = mod_4529_bufferize.operation;
    Operation_IFC mod_4529 <- mkDebugOperation(mod_4529_inner, "mod_4529");
    PMU_IFC mod_4530_bufferize <- mkPMU(2);
    Operation_IFC mod_4530_inner = mod_4530_bufferize.operation;
    Operation_IFC mod_4530 <- mkDebugOperation(mod_4530_inner, "mod_4530");
    Operation_IFC mod_4531_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4531 <- mkDebugOperation(mod_4531_inner, "mod_4531");
    Operation_IFC mod_4532_inner <- mkFlatten(1);
    Operation_IFC mod_4532 <- mkDebugOperation(mod_4532_inner, "mod_4532");
    Operation_IFC mod_4533_inner <- mkFlatten(0);
    Operation_IFC mod_4533 <- mkDebugOperation(mod_4533_inner, "mod_4533");
    Operation_IFC mod_4534_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4534 <- mkDebugOperation(mod_4534_inner, "mod_4534");
    Operation_IFC mod_4535_inner <- mkUnaryMap(1686, silu_tile);
    Operation_IFC mod_4535 <- mkDebugOperation(mod_4535_inner, "mod_4535");
    Operation_IFC mod_4536_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4536 <- mkDebugOperation(mod_4536_inner, "mod_4536");
    Operation_IFC mod_4537_inner <- mkBinaryMap(1558, matmul_t_tile);
    Operation_IFC mod_4537 <- mkDebugOperation(mod_4537_inner, "mod_4537");
    PMU_IFC mod_4538_bufferize <- mkPMU(2);
    Operation_IFC mod_4538_inner = mod_4538_bufferize.operation;
    Operation_IFC mod_4538 <- mkDebugOperation(mod_4538_inner, "mod_4538");
    Operation_IFC mod_4539_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4539 <- mkDebugOperation(mod_4539_inner, "mod_4539");
    Operation_IFC mod_4540_inner <- mkFlatten(1);
    Operation_IFC mod_4540 <- mkDebugOperation(mod_4540_inner, "mod_4540");
    Operation_IFC mod_4541_inner <- mkFlatten(0);
    Operation_IFC mod_4541 <- mkDebugOperation(mod_4541_inner, "mod_4541");
    PMU_IFC mod_4542_bufferize <- mkPMU(1);
    Operation_IFC mod_4542_inner = mod_4542_bufferize.operation;
    Operation_IFC mod_4542 <- mkDebugOperation(mod_4542_inner, "mod_4542");
    Operation_IFC mod_4543_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4543 <- mkDebugOperation(mod_4543_inner, "mod_4543");
    PMU_IFC mod_4544_bufferize <- mkPMU(2);
    Operation_IFC mod_4544_inner = mod_4544_bufferize.operation;
    Operation_IFC mod_4544 <- mkDebugOperation(mod_4544_inner, "mod_4544");
    Operation_IFC mod_4545_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4545 <- mkDebugOperation(mod_4545_inner, "mod_4545");
    Operation_IFC mod_4546_inner <- mkFlatten(1);
    Operation_IFC mod_4546 <- mkDebugOperation(mod_4546_inner, "mod_4546");
    Operation_IFC mod_4547_inner <- mkFlatten(0);
    Operation_IFC mod_4547 <- mkDebugOperation(mod_4547_inner, "mod_4547");
    Operation_IFC mod_4548_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4548 <- mkDebugOperation(mod_4548_inner, "mod_4548");
    Operation_IFC mod_4549_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4549 <- mkDebugOperation(mod_4549_inner, "mod_4549");
    PMU_IFC mod_4550_bufferize <- mkPMU(2);
    Operation_IFC mod_4550_inner = mod_4550_bufferize.operation;
    Operation_IFC mod_4550 <- mkDebugOperation(mod_4550_inner, "mod_4550");
    rule rule_5831;
        ChannelMessage t;
        t <- mod_4529.get(0);
        mod_4529.put(1, t);
    endrule
    rule rule_5832;
        ChannelMessage t;
        t <- mod_4541.get(0);
        mod_4540.put(0, t);
    endrule
    rule rule_5833;
        ChannelMessage t;
        t <- mod_4534.get(0);
        mod_4522.put(1, t);
    endrule
    rule rule_5834;
        ChannelMessage t;
        t <- mod_4519.get(0);
        mod_4520.put(0, t);
    endrule
    rule rule_5835;
        ChannelMessage t;
        t <- mod_4542.get(0);
        mod_4543.put(0, t);
    endrule
    rule rule_5836;
        ChannelMessage t;
        t <- mod_4516.get(1);
        mod_4517.put(0, t);
    endrule
    rule rule_5837;
        ChannelMessage t;
        t <- mod_4530.get(0);
        mod_4531.put(0, t);
    endrule
    rule rule_5838;
        ChannelMessage t;
        t <- mod_4512.get(0);
        mod_4513.put(0, t);
    endrule
    rule rule_5839;
        ChannelMessage t;
        t <- mod_4545.get(0);
        mod_4544.put(1, t);
    endrule
    rule rule_5840;
        ChannelMessage t;
        t <- mod_4521.get(0);
        mod_4522.put(0, t);
    endrule
    rule rule_5841;
        ChannelMessage t;
        t <- mod_4518.get(1);
        mod_4519.put(0, t);
    endrule
    rule rule_5842;
        ChannelMessage t;
        t <- mod_4515.get(3);
        mod_4516.put(0, t);
    endrule
    rule rule_5843;
        ChannelMessage t;
        t <- mod_4517.get(0);
        mod_4542.put(0, t);
    endrule
    rule rule_5844;
        ChannelMessage t;
        t <- mod_4524.get(0);
        mod_4525.put(0, t);
    endrule
    rule rule_5845;
        ChannelMessage t;
        t <- mod_4538.get(1);
        mod_4537.put(1, t);
    endrule
    rule rule_5846;
        ChannelMessage t;
        t <- mod_4543.get(0);
        mod_4542.put(1, t);
    endrule
    rule rule_5847;
        ChannelMessage t;
        t <- mod_4536.get(0);
        mod_4535.put(0, t);
    endrule
    rule rule_5848;
        ChannelMessage t;
        t <- mod_4550.get(0);
        mod_4550.put(1, t);
    endrule
    rule rule_5849;
        ChannelMessage t;
        t <- mod_4523.get(0);
        mod_4524.put(0, t);
    endrule
    rule rule_5850;
        ChannelMessage t;
        t <- mod_4520.get(0);
        mod_4521.put(0, t);
    endrule
    rule rule_5851;
        ChannelMessage t;
        t <- mod_4526.get(0);
        mod_4528.put(0, t);
    endrule
    rule rule_5852;
        ChannelMessage t;
        t <- mod_4528.get(1);
        mod_4526.put(1, t);
    endrule
    rule rule_5853;
        ChannelMessage t;
        t <- mod_4526.get(1);
        mod_4527.put(1, t);
    endrule
    rule rule_5854;
        ChannelMessage t;
        t <- mod_4533.get(0);
        mod_4532.put(0, t);
    endrule
    rule rule_5855;
        ChannelMessage t;
        t <- mod_4522.get(1);
        mod_4523.put(0, t);
    endrule
    rule rule_5856;
        ChannelMessage t;
        t <- mod_4532.get(0);
        mod_4530.put(0, t);
    endrule
    rule rule_5857;
        ChannelMessage t;
        t <- mod_4544.get(1);
        mod_4519.put(1, t);
    endrule
    rule rule_5858;
        ChannelMessage t;
        t <- mod_4522.get(0);
        mod_4534.put(0, t);
    endrule
    rule rule_5859;
        ChannelMessage t;
        t <- mod_4547.get(0);
        mod_4546.put(0, t);
    endrule
    rule rule_5860;
        ChannelMessage t;
        t <- mod_4517.get(1);
        mod_4518.put(0, t);
    endrule
    rule rule_5861;
        ChannelMessage t;
        t <- mod_4514.get(1);
        mod_4515.put(0, t);
    endrule
    rule rule_5862;
        ChannelMessage t;
        t <- mod_4529.get(1);
        mod_4525.put(1, t);
    endrule
    rule rule_5863;
        ChannelMessage t;
        t <- mod_4544.get(0);
        mod_4545.put(0, t);
    endrule
    rule rule_5864;
        ChannelMessage t;
        t <- mod_4528.get(0);
        mod_4528.put(1, t);
    endrule
    rule rule_5865;
        ChannelMessage t;
        t <- mod_4530.get(1);
        mod_4523.put(1, t);
    endrule
    rule rule_5866;
        ChannelMessage t;
        t <- mod_4542.get(1);
        mod_4537.put(0, t);
    endrule
    rule rule_5867;
        ChannelMessage t;
        t <- mod_4518.get(0);
        mod_4548.put(0, t);
    endrule
    rule rule_5868;
        ChannelMessage t;
        t <- mod_4525.get(0);
        mod_4529.put(0, t);
    endrule
    rule rule_5869;
        ChannelMessage t;
        t <- mod_4548.get(0);
        mod_4518.put(1, t);
    endrule
    rule rule_5870;
        ChannelMessage t;
        t <- mod_4546.get(0);
        mod_4544.put(0, t);
    endrule
    rule rule_5871;
        ChannelMessage t;
        t <- mod_4550.get(1);
        mod_4514.put(1, t);
    endrule
    rule rule_5872;
        ChannelMessage t;
        t <- mod_4525.get(1);
        mod_4526.put(0, t);
    endrule
    rule rule_5873;
        ChannelMessage t;
        t <- mod_4535.get(0);
        mod_4521.put(1, t);
    endrule
    rule rule_5874;
        ChannelMessage t;
        t <- mod_4531.get(0);
        mod_4530.put(1, t);
    endrule
    rule rule_5875;
        ChannelMessage t;
        t <- mod_4539.get(0);
        mod_4538.put(1, t);
    endrule
    rule rule_5876;
        ChannelMessage t;
        t <- mod_4513.get(0);
        mod_4514.put(0, t);
    endrule
    rule rule_5877;
        ChannelMessage t;
        t <- mod_4537.get(0);
        mod_4536.put(0, t);
    endrule
    rule rule_5878;
        ChannelMessage t;
        t <- mod_4514.get(0);
        mod_4550.put(0, t);
    endrule
    rule rule_5879;
        ChannelMessage t;
        t <- mod_4511.get(0);
        mod_4512.put(0, t);
    endrule
    rule rule_5880;
        ChannelMessage t;
        t <- mod_4540.get(0);
        mod_4538.put(0, t);
    endrule
    rule rule_5881;
        ChannelMessage t;
        t <- mod_4549.get(0);
        mod_4516.put(1, t);
    endrule
    rule rule_5882;
        ChannelMessage t;
        t <- mod_4516.get(0);
        mod_4549.put(0, t);
    endrule
    rule rule_5883;
        ChannelMessage t;
        t <- mod_4538.get(0);
        mod_4539.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4511.put(0, t);
        end
        if (i == 1) begin
            mod_4527.put(0, t);
        end
        if (i == 2) begin
            mod_4533.put(0, t);
        end
        if (i == 3) begin
            mod_4541.put(0, t);
        end
        if (i == 4) begin
            mod_4547.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_4515.get(0);
        end
        if (i == 2) begin
            t <- mod_4515.get(1);
        end
        if (i == 0) begin
            t <- mod_4515.get(2);
        end
        if (i == 1) begin
            t <- mod_4527.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6145 (Operation_IFC);
    Operation_IFC mod_4552_inner <- mkReshape(2, 64);
    Operation_IFC mod_4552 <- mkDebugOperation(mod_4552_inner, "mod_4552");
    Operation_IFC mod_4553_inner <- mkFlatten(1);
    Operation_IFC mod_4553 <- mkDebugOperation(mod_4553_inner, "mod_4553");
    Operation_IFC mod_4554_inner <- mkFlatten(2);
    Operation_IFC mod_4554 <- mkDebugOperation(mod_4554_inner, "mod_4554");
    Operation_IFC mod_4555_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4555 <- mkDebugOperation(mod_4555_inner, "mod_4555");
    Broadcast_IFC#(4) mod_4556_inner <- mkBroadcast(4);
    Operation_IFC mod_4556 <- mkDebugOperation(mod_4556_inner.op, "mod_4556");
    PMU_IFC mod_4557_bufferize <- mkPMU(2);
    Operation_IFC mod_4557_inner = mod_4557_bufferize.operation;
    Operation_IFC mod_4557 <- mkDebugOperation(mod_4557_inner, "mod_4557");
    Broadcast_IFC#(2) mod_4558_inner <- mkBroadcast(2);
    Operation_IFC mod_4558 <- mkDebugOperation(mod_4558_inner.op, "mod_4558");
    PMU_IFC mod_4559_bufferize <- mkPMU(1);
    Operation_IFC mod_4559_inner = mod_4559_bufferize.operation;
    Operation_IFC mod_4559 <- mkDebugOperation(mod_4559_inner, "mod_4559");
    Operation_IFC mod_4560_inner <- mkBinaryMap(1045, matmul_t_tile);
    Operation_IFC mod_4560 <- mkDebugOperation(mod_4560_inner, "mod_4560");
    Operation_IFC mod_4561_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4561 <- mkDebugOperation(mod_4561_inner, "mod_4561");
    Operation_IFC mod_4562_inner <- mkBinaryMap(1813, mul_tile);
    Operation_IFC mod_4562 <- mkDebugOperation(mod_4562_inner, "mod_4562");
    PMU_IFC mod_4563_bufferize <- mkPMU(1);
    Operation_IFC mod_4563_inner = mod_4563_bufferize.operation;
    Operation_IFC mod_4563 <- mkDebugOperation(mod_4563_inner, "mod_4563");
    Operation_IFC mod_4564_inner <- mkBinaryMap(2341, matmul_t_tile);
    Operation_IFC mod_4564 <- mkDebugOperation(mod_4564_inner, "mod_4564");
    Operation_IFC mod_4565_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4565 <- mkDebugOperation(mod_4565_inner, "mod_4565");
    Operation_IFC mod_4566_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4566 <- mkDebugOperation(mod_4566_inner, "mod_4566");
    Operation_IFC mod_4567_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4567 <- mkDebugOperation(mod_4567_inner, "mod_4567");
    Operation_IFC mod_4568_inner <- mkBinaryMap(2712, mul_tile);
    Operation_IFC mod_4568 <- mkDebugOperation(mod_4568_inner, "mod_4568");
    PMU_IFC mod_4569_bufferize <- mkPMU(1);
    Operation_IFC mod_4569_inner = mod_4569_bufferize.operation;
    Operation_IFC mod_4569 <- mkDebugOperation(mod_4569_inner, "mod_4569");
    PMU_IFC mod_4570_bufferize <- mkPMU(2);
    Operation_IFC mod_4570_inner = mod_4570_bufferize.operation;
    Operation_IFC mod_4570 <- mkDebugOperation(mod_4570_inner, "mod_4570");
    PMU_IFC mod_4571_bufferize <- mkPMU(2);
    Operation_IFC mod_4571_inner = mod_4571_bufferize.operation;
    Operation_IFC mod_4571 <- mkDebugOperation(mod_4571_inner, "mod_4571");
    Operation_IFC mod_4572_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4572 <- mkDebugOperation(mod_4572_inner, "mod_4572");
    Operation_IFC mod_4573_inner <- mkFlatten(1);
    Operation_IFC mod_4573 <- mkDebugOperation(mod_4573_inner, "mod_4573");
    Operation_IFC mod_4574_inner <- mkFlatten(0);
    Operation_IFC mod_4574 <- mkDebugOperation(mod_4574_inner, "mod_4574");
    Operation_IFC mod_4575_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4575 <- mkDebugOperation(mod_4575_inner, "mod_4575");
    Operation_IFC mod_4576_inner <- mkUnaryMap(1685, silu_tile);
    Operation_IFC mod_4576 <- mkDebugOperation(mod_4576_inner, "mod_4576");
    Operation_IFC mod_4577_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4577 <- mkDebugOperation(mod_4577_inner, "mod_4577");
    Operation_IFC mod_4578_inner <- mkBinaryMap(1557, matmul_t_tile);
    Operation_IFC mod_4578 <- mkDebugOperation(mod_4578_inner, "mod_4578");
    PMU_IFC mod_4579_bufferize <- mkPMU(2);
    Operation_IFC mod_4579_inner = mod_4579_bufferize.operation;
    Operation_IFC mod_4579 <- mkDebugOperation(mod_4579_inner, "mod_4579");
    Operation_IFC mod_4580_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4580 <- mkDebugOperation(mod_4580_inner, "mod_4580");
    Operation_IFC mod_4581_inner <- mkFlatten(1);
    Operation_IFC mod_4581 <- mkDebugOperation(mod_4581_inner, "mod_4581");
    Operation_IFC mod_4582_inner <- mkFlatten(0);
    Operation_IFC mod_4582 <- mkDebugOperation(mod_4582_inner, "mod_4582");
    PMU_IFC mod_4583_bufferize <- mkPMU(1);
    Operation_IFC mod_4583_inner = mod_4583_bufferize.operation;
    Operation_IFC mod_4583 <- mkDebugOperation(mod_4583_inner, "mod_4583");
    Operation_IFC mod_4584_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4584 <- mkDebugOperation(mod_4584_inner, "mod_4584");
    PMU_IFC mod_4585_bufferize <- mkPMU(2);
    Operation_IFC mod_4585_inner = mod_4585_bufferize.operation;
    Operation_IFC mod_4585 <- mkDebugOperation(mod_4585_inner, "mod_4585");
    Operation_IFC mod_4586_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4586 <- mkDebugOperation(mod_4586_inner, "mod_4586");
    Operation_IFC mod_4587_inner <- mkFlatten(1);
    Operation_IFC mod_4587 <- mkDebugOperation(mod_4587_inner, "mod_4587");
    Operation_IFC mod_4588_inner <- mkFlatten(0);
    Operation_IFC mod_4588 <- mkDebugOperation(mod_4588_inner, "mod_4588");
    Operation_IFC mod_4589_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4589 <- mkDebugOperation(mod_4589_inner, "mod_4589");
    Operation_IFC mod_4590_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4590 <- mkDebugOperation(mod_4590_inner, "mod_4590");
    PMU_IFC mod_4591_bufferize <- mkPMU(2);
    Operation_IFC mod_4591_inner = mod_4591_bufferize.operation;
    Operation_IFC mod_4591 <- mkDebugOperation(mod_4591_inner, "mod_4591");
    rule rule_5884;
        ChannelMessage t;
        t <- mod_4588.get(0);
        mod_4587.put(0, t);
    endrule
    rule rule_5885;
        ChannelMessage t;
        t <- mod_4577.get(0);
        mod_4576.put(0, t);
    endrule
    rule rule_5886;
        ChannelMessage t;
        t <- mod_4558.get(0);
        mod_4583.put(0, t);
    endrule
    rule rule_5887;
        ChannelMessage t;
        t <- mod_4587.get(0);
        mod_4585.put(0, t);
    endrule
    rule rule_5888;
        ChannelMessage t;
        t <- mod_4567.get(0);
        mod_4569.put(0, t);
    endrule
    rule rule_5889;
        ChannelMessage t;
        t <- mod_4565.get(0);
        mod_4566.put(0, t);
    endrule
    rule rule_5890;
        ChannelMessage t;
        t <- mod_4566.get(1);
        mod_4567.put(0, t);
    endrule
    rule rule_5891;
        ChannelMessage t;
        t <- mod_4564.get(0);
        mod_4565.put(0, t);
    endrule
    rule rule_5892;
        ChannelMessage t;
        t <- mod_4571.get(0);
        mod_4572.put(0, t);
    endrule
    rule rule_5893;
        ChannelMessage t;
        t <- mod_4579.get(1);
        mod_4578.put(1, t);
    endrule
    rule rule_5894;
        ChannelMessage t;
        t <- mod_4584.get(0);
        mod_4583.put(1, t);
    endrule
    rule rule_5895;
        ChannelMessage t;
        t <- mod_4563.get(1);
        mod_4564.put(0, t);
    endrule
    rule rule_5896;
        ChannelMessage t;
        t <- mod_4563.get(0);
        mod_4575.put(0, t);
    endrule
    rule rule_5897;
        ChannelMessage t;
        t <- mod_4578.get(0);
        mod_4577.put(0, t);
    endrule
    rule rule_5898;
        ChannelMessage t;
        t <- mod_4585.get(0);
        mod_4586.put(0, t);
    endrule
    rule rule_5899;
        ChannelMessage t;
        t <- mod_4574.get(0);
        mod_4573.put(0, t);
    endrule
    rule rule_5900;
        ChannelMessage t;
        t <- mod_4562.get(0);
        mod_4563.put(0, t);
    endrule
    rule rule_5901;
        ChannelMessage t;
        t <- mod_4579.get(0);
        mod_4580.put(0, t);
    endrule
    rule rule_5902;
        ChannelMessage t;
        t <- mod_4555.get(1);
        mod_4556.put(0, t);
    endrule
    rule rule_5903;
        ChannelMessage t;
        t <- mod_4583.get(1);
        mod_4578.put(0, t);
    endrule
    rule rule_5904;
        ChannelMessage t;
        t <- mod_4591.get(1);
        mod_4555.put(1, t);
    endrule
    rule rule_5905;
        ChannelMessage t;
        t <- mod_4570.get(0);
        mod_4570.put(1, t);
    endrule
    rule rule_5906;
        ChannelMessage t;
        t <- mod_4573.get(0);
        mod_4571.put(0, t);
    endrule
    rule rule_5907;
        ChannelMessage t;
        t <- mod_4580.get(0);
        mod_4579.put(1, t);
    endrule
    rule rule_5908;
        ChannelMessage t;
        t <- mod_4583.get(0);
        mod_4584.put(0, t);
    endrule
    rule rule_5909;
        ChannelMessage t;
        t <- mod_4585.get(1);
        mod_4560.put(1, t);
    endrule
    rule rule_5910;
        ChannelMessage t;
        t <- mod_4555.get(0);
        mod_4591.put(0, t);
    endrule
    rule rule_5911;
        ChannelMessage t;
        t <- mod_4591.get(0);
        mod_4591.put(1, t);
    endrule
    rule rule_5912;
        ChannelMessage t;
        t <- mod_4566.get(0);
        mod_4570.put(0, t);
    endrule
    rule rule_5913;
        ChannelMessage t;
        t <- mod_4586.get(0);
        mod_4585.put(1, t);
    endrule
    rule rule_5914;
        ChannelMessage t;
        t <- mod_4567.get(1);
        mod_4568.put(1, t);
    endrule
    rule rule_5915;
        ChannelMessage t;
        t <- mod_4572.get(0);
        mod_4571.put(1, t);
    endrule
    rule rule_5916;
        ChannelMessage t;
        t <- mod_4581.get(0);
        mod_4579.put(0, t);
    endrule
    rule rule_5917;
        ChannelMessage t;
        t <- mod_4557.get(0);
        mod_4590.put(0, t);
    endrule
    rule rule_5918;
        ChannelMessage t;
        t <- mod_4552.get(0);
        mod_4553.put(0, t);
    endrule
    rule rule_5919;
        ChannelMessage t;
        t <- mod_4582.get(0);
        mod_4581.put(0, t);
    endrule
    rule rule_5920;
        ChannelMessage t;
        t <- mod_4569.get(1);
        mod_4567.put(1, t);
    endrule
    rule rule_5921;
        ChannelMessage t;
        t <- mod_4553.get(0);
        mod_4554.put(0, t);
    endrule
    rule rule_5922;
        ChannelMessage t;
        t <- mod_4559.get(0);
        mod_4589.put(0, t);
    endrule
    rule rule_5923;
        ChannelMessage t;
        t <- mod_4559.get(1);
        mod_4560.put(0, t);
    endrule
    rule rule_5924;
        ChannelMessage t;
        t <- mod_4556.get(3);
        mod_4557.put(0, t);
    endrule
    rule rule_5925;
        ChannelMessage t;
        t <- mod_4576.get(0);
        mod_4562.put(1, t);
    endrule
    rule rule_5926;
        ChannelMessage t;
        t <- mod_4570.get(1);
        mod_4566.put(1, t);
    endrule
    rule rule_5927;
        ChannelMessage t;
        t <- mod_4590.get(0);
        mod_4557.put(1, t);
    endrule
    rule rule_5928;
        ChannelMessage t;
        t <- mod_4560.get(0);
        mod_4561.put(0, t);
    endrule
    rule rule_5929;
        ChannelMessage t;
        t <- mod_4569.get(0);
        mod_4569.put(1, t);
    endrule
    rule rule_5930;
        ChannelMessage t;
        t <- mod_4561.get(0);
        mod_4562.put(0, t);
    endrule
    rule rule_5931;
        ChannelMessage t;
        t <- mod_4558.get(1);
        mod_4559.put(0, t);
    endrule
    rule rule_5932;
        ChannelMessage t;
        t <- mod_4557.get(1);
        mod_4558.put(0, t);
    endrule
    rule rule_5933;
        ChannelMessage t;
        t <- mod_4571.get(1);
        mod_4564.put(1, t);
    endrule
    rule rule_5934;
        ChannelMessage t;
        t <- mod_4554.get(0);
        mod_4555.put(0, t);
    endrule
    rule rule_5935;
        ChannelMessage t;
        t <- mod_4575.get(0);
        mod_4563.put(1, t);
    endrule
    rule rule_5936;
        ChannelMessage t;
        t <- mod_4589.get(0);
        mod_4559.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4552.put(0, t);
        end
        if (i == 1) begin
            mod_4568.put(0, t);
        end
        if (i == 2) begin
            mod_4574.put(0, t);
        end
        if (i == 3) begin
            mod_4582.put(0, t);
        end
        if (i == 4) begin
            mod_4588.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_4556.get(0);
        end
        if (i == 0) begin
            t <- mod_4556.get(1);
        end
        if (i == 2) begin
            t <- mod_4556.get(2);
        end
        if (i == 3) begin
            t <- mod_4568.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6146 (Operation_IFC);
    Operation_IFC mod_4593_inner <- mkReshape(2, 64);
    Operation_IFC mod_4593 <- mkDebugOperation(mod_4593_inner, "mod_4593");
    Operation_IFC mod_4594_inner <- mkFlatten(1);
    Operation_IFC mod_4594 <- mkDebugOperation(mod_4594_inner, "mod_4594");
    Operation_IFC mod_4595_inner <- mkFlatten(2);
    Operation_IFC mod_4595 <- mkDebugOperation(mod_4595_inner, "mod_4595");
    Operation_IFC mod_4596_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4596 <- mkDebugOperation(mod_4596_inner, "mod_4596");
    Broadcast_IFC#(4) mod_4597_inner <- mkBroadcast(4);
    Operation_IFC mod_4597 <- mkDebugOperation(mod_4597_inner.op, "mod_4597");
    PMU_IFC mod_4598_bufferize <- mkPMU(2);
    Operation_IFC mod_4598_inner = mod_4598_bufferize.operation;
    Operation_IFC mod_4598 <- mkDebugOperation(mod_4598_inner, "mod_4598");
    Broadcast_IFC#(2) mod_4599_inner <- mkBroadcast(2);
    Operation_IFC mod_4599 <- mkDebugOperation(mod_4599_inner.op, "mod_4599");
    PMU_IFC mod_4600_bufferize <- mkPMU(1);
    Operation_IFC mod_4600_inner = mod_4600_bufferize.operation;
    Operation_IFC mod_4600 <- mkDebugOperation(mod_4600_inner, "mod_4600");
    Operation_IFC mod_4601_inner <- mkBinaryMap(1044, matmul_t_tile);
    Operation_IFC mod_4601 <- mkDebugOperation(mod_4601_inner, "mod_4601");
    Operation_IFC mod_4602_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4602 <- mkDebugOperation(mod_4602_inner, "mod_4602");
    Operation_IFC mod_4603_inner <- mkBinaryMap(1812, mul_tile);
    Operation_IFC mod_4603 <- mkDebugOperation(mod_4603_inner, "mod_4603");
    PMU_IFC mod_4604_bufferize <- mkPMU(1);
    Operation_IFC mod_4604_inner = mod_4604_bufferize.operation;
    Operation_IFC mod_4604 <- mkDebugOperation(mod_4604_inner, "mod_4604");
    Operation_IFC mod_4605_inner <- mkBinaryMap(2339, matmul_t_tile);
    Operation_IFC mod_4605 <- mkDebugOperation(mod_4605_inner, "mod_4605");
    Operation_IFC mod_4606_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4606 <- mkDebugOperation(mod_4606_inner, "mod_4606");
    Operation_IFC mod_4607_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4607 <- mkDebugOperation(mod_4607_inner, "mod_4607");
    Operation_IFC mod_4608_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4608 <- mkDebugOperation(mod_4608_inner, "mod_4608");
    Operation_IFC mod_4609_inner <- mkBinaryMap(2711, mul_tile);
    Operation_IFC mod_4609 <- mkDebugOperation(mod_4609_inner, "mod_4609");
    PMU_IFC mod_4610_bufferize <- mkPMU(1);
    Operation_IFC mod_4610_inner = mod_4610_bufferize.operation;
    Operation_IFC mod_4610 <- mkDebugOperation(mod_4610_inner, "mod_4610");
    PMU_IFC mod_4611_bufferize <- mkPMU(2);
    Operation_IFC mod_4611_inner = mod_4611_bufferize.operation;
    Operation_IFC mod_4611 <- mkDebugOperation(mod_4611_inner, "mod_4611");
    PMU_IFC mod_4612_bufferize <- mkPMU(2);
    Operation_IFC mod_4612_inner = mod_4612_bufferize.operation;
    Operation_IFC mod_4612 <- mkDebugOperation(mod_4612_inner, "mod_4612");
    Operation_IFC mod_4613_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4613 <- mkDebugOperation(mod_4613_inner, "mod_4613");
    Operation_IFC mod_4614_inner <- mkFlatten(1);
    Operation_IFC mod_4614 <- mkDebugOperation(mod_4614_inner, "mod_4614");
    Operation_IFC mod_4615_inner <- mkFlatten(0);
    Operation_IFC mod_4615 <- mkDebugOperation(mod_4615_inner, "mod_4615");
    Operation_IFC mod_4616_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4616 <- mkDebugOperation(mod_4616_inner, "mod_4616");
    Operation_IFC mod_4617_inner <- mkUnaryMap(1684, silu_tile);
    Operation_IFC mod_4617 <- mkDebugOperation(mod_4617_inner, "mod_4617");
    Operation_IFC mod_4618_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4618 <- mkDebugOperation(mod_4618_inner, "mod_4618");
    Operation_IFC mod_4619_inner <- mkBinaryMap(1556, matmul_t_tile);
    Operation_IFC mod_4619 <- mkDebugOperation(mod_4619_inner, "mod_4619");
    PMU_IFC mod_4620_bufferize <- mkPMU(2);
    Operation_IFC mod_4620_inner = mod_4620_bufferize.operation;
    Operation_IFC mod_4620 <- mkDebugOperation(mod_4620_inner, "mod_4620");
    Operation_IFC mod_4621_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4621 <- mkDebugOperation(mod_4621_inner, "mod_4621");
    Operation_IFC mod_4622_inner <- mkFlatten(1);
    Operation_IFC mod_4622 <- mkDebugOperation(mod_4622_inner, "mod_4622");
    Operation_IFC mod_4623_inner <- mkFlatten(0);
    Operation_IFC mod_4623 <- mkDebugOperation(mod_4623_inner, "mod_4623");
    PMU_IFC mod_4624_bufferize <- mkPMU(1);
    Operation_IFC mod_4624_inner = mod_4624_bufferize.operation;
    Operation_IFC mod_4624 <- mkDebugOperation(mod_4624_inner, "mod_4624");
    Operation_IFC mod_4625_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4625 <- mkDebugOperation(mod_4625_inner, "mod_4625");
    PMU_IFC mod_4626_bufferize <- mkPMU(2);
    Operation_IFC mod_4626_inner = mod_4626_bufferize.operation;
    Operation_IFC mod_4626 <- mkDebugOperation(mod_4626_inner, "mod_4626");
    Operation_IFC mod_4627_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4627 <- mkDebugOperation(mod_4627_inner, "mod_4627");
    Operation_IFC mod_4628_inner <- mkFlatten(1);
    Operation_IFC mod_4628 <- mkDebugOperation(mod_4628_inner, "mod_4628");
    Operation_IFC mod_4629_inner <- mkFlatten(0);
    Operation_IFC mod_4629 <- mkDebugOperation(mod_4629_inner, "mod_4629");
    Operation_IFC mod_4630_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4630 <- mkDebugOperation(mod_4630_inner, "mod_4630");
    Operation_IFC mod_4631_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4631 <- mkDebugOperation(mod_4631_inner, "mod_4631");
    PMU_IFC mod_4632_bufferize <- mkPMU(2);
    Operation_IFC mod_4632_inner = mod_4632_bufferize.operation;
    Operation_IFC mod_4632 <- mkDebugOperation(mod_4632_inner, "mod_4632");
    rule rule_5937;
        ChannelMessage t;
        t <- mod_4602.get(0);
        mod_4603.put(0, t);
    endrule
    rule rule_5938;
        ChannelMessage t;
        t <- mod_4596.get(0);
        mod_4632.put(0, t);
    endrule
    rule rule_5939;
        ChannelMessage t;
        t <- mod_4611.get(1);
        mod_4607.put(1, t);
    endrule
    rule rule_5940;
        ChannelMessage t;
        t <- mod_4614.get(0);
        mod_4612.put(0, t);
    endrule
    rule rule_5941;
        ChannelMessage t;
        t <- mod_4604.get(0);
        mod_4616.put(0, t);
    endrule
    rule rule_5942;
        ChannelMessage t;
        t <- mod_4599.get(0);
        mod_4624.put(0, t);
    endrule
    rule rule_5943;
        ChannelMessage t;
        t <- mod_4616.get(0);
        mod_4604.put(1, t);
    endrule
    rule rule_5944;
        ChannelMessage t;
        t <- mod_4603.get(0);
        mod_4604.put(0, t);
    endrule
    rule rule_5945;
        ChannelMessage t;
        t <- mod_4593.get(0);
        mod_4594.put(0, t);
    endrule
    rule rule_5946;
        ChannelMessage t;
        t <- mod_4624.get(1);
        mod_4619.put(0, t);
    endrule
    rule rule_5947;
        ChannelMessage t;
        t <- mod_4604.get(1);
        mod_4605.put(0, t);
    endrule
    rule rule_5948;
        ChannelMessage t;
        t <- mod_4632.get(1);
        mod_4596.put(1, t);
    endrule
    rule rule_5949;
        ChannelMessage t;
        t <- mod_4620.get(0);
        mod_4621.put(0, t);
    endrule
    rule rule_5950;
        ChannelMessage t;
        t <- mod_4629.get(0);
        mod_4628.put(0, t);
    endrule
    rule rule_5951;
        ChannelMessage t;
        t <- mod_4631.get(0);
        mod_4598.put(1, t);
    endrule
    rule rule_5952;
        ChannelMessage t;
        t <- mod_4618.get(0);
        mod_4617.put(0, t);
    endrule
    rule rule_5953;
        ChannelMessage t;
        t <- mod_4607.get(1);
        mod_4608.put(0, t);
    endrule
    rule rule_5954;
        ChannelMessage t;
        t <- mod_4598.get(0);
        mod_4631.put(0, t);
    endrule
    rule rule_5955;
        ChannelMessage t;
        t <- mod_4628.get(0);
        mod_4626.put(0, t);
    endrule
    rule rule_5956;
        ChannelMessage t;
        t <- mod_4598.get(1);
        mod_4599.put(0, t);
    endrule
    rule rule_5957;
        ChannelMessage t;
        t <- mod_4619.get(0);
        mod_4618.put(0, t);
    endrule
    rule rule_5958;
        ChannelMessage t;
        t <- mod_4611.get(0);
        mod_4611.put(1, t);
    endrule
    rule rule_5959;
        ChannelMessage t;
        t <- mod_4621.get(0);
        mod_4620.put(1, t);
    endrule
    rule rule_5960;
        ChannelMessage t;
        t <- mod_4610.get(0);
        mod_4610.put(1, t);
    endrule
    rule rule_5961;
        ChannelMessage t;
        t <- mod_4625.get(0);
        mod_4624.put(1, t);
    endrule
    rule rule_5962;
        ChannelMessage t;
        t <- mod_4596.get(1);
        mod_4597.put(0, t);
    endrule
    rule rule_5963;
        ChannelMessage t;
        t <- mod_4599.get(1);
        mod_4600.put(0, t);
    endrule
    rule rule_5964;
        ChannelMessage t;
        t <- mod_4607.get(0);
        mod_4611.put(0, t);
    endrule
    rule rule_5965;
        ChannelMessage t;
        t <- mod_4620.get(1);
        mod_4619.put(1, t);
    endrule
    rule rule_5966;
        ChannelMessage t;
        t <- mod_4600.get(1);
        mod_4601.put(0, t);
    endrule
    rule rule_5967;
        ChannelMessage t;
        t <- mod_4623.get(0);
        mod_4622.put(0, t);
    endrule
    rule rule_5968;
        ChannelMessage t;
        t <- mod_4610.get(1);
        mod_4608.put(1, t);
    endrule
    rule rule_5969;
        ChannelMessage t;
        t <- mod_4626.get(1);
        mod_4601.put(1, t);
    endrule
    rule rule_5970;
        ChannelMessage t;
        t <- mod_4622.get(0);
        mod_4620.put(0, t);
    endrule
    rule rule_5971;
        ChannelMessage t;
        t <- mod_4605.get(0);
        mod_4606.put(0, t);
    endrule
    rule rule_5972;
        ChannelMessage t;
        t <- mod_4597.get(3);
        mod_4598.put(0, t);
    endrule
    rule rule_5973;
        ChannelMessage t;
        t <- mod_4608.get(1);
        mod_4609.put(1, t);
    endrule
    rule rule_5974;
        ChannelMessage t;
        t <- mod_4601.get(0);
        mod_4602.put(0, t);
    endrule
    rule rule_5975;
        ChannelMessage t;
        t <- mod_4608.get(0);
        mod_4610.put(0, t);
    endrule
    rule rule_5976;
        ChannelMessage t;
        t <- mod_4624.get(0);
        mod_4625.put(0, t);
    endrule
    rule rule_5977;
        ChannelMessage t;
        t <- mod_4630.get(0);
        mod_4600.put(1, t);
    endrule
    rule rule_5978;
        ChannelMessage t;
        t <- mod_4612.get(1);
        mod_4605.put(1, t);
    endrule
    rule rule_5979;
        ChannelMessage t;
        t <- mod_4594.get(0);
        mod_4595.put(0, t);
    endrule
    rule rule_5980;
        ChannelMessage t;
        t <- mod_4613.get(0);
        mod_4612.put(1, t);
    endrule
    rule rule_5981;
        ChannelMessage t;
        t <- mod_4627.get(0);
        mod_4626.put(1, t);
    endrule
    rule rule_5982;
        ChannelMessage t;
        t <- mod_4632.get(0);
        mod_4632.put(1, t);
    endrule
    rule rule_5983;
        ChannelMessage t;
        t <- mod_4615.get(0);
        mod_4614.put(0, t);
    endrule
    rule rule_5984;
        ChannelMessage t;
        t <- mod_4606.get(0);
        mod_4607.put(0, t);
    endrule
    rule rule_5985;
        ChannelMessage t;
        t <- mod_4612.get(0);
        mod_4613.put(0, t);
    endrule
    rule rule_5986;
        ChannelMessage t;
        t <- mod_4617.get(0);
        mod_4603.put(1, t);
    endrule
    rule rule_5987;
        ChannelMessage t;
        t <- mod_4600.get(0);
        mod_4630.put(0, t);
    endrule
    rule rule_5988;
        ChannelMessage t;
        t <- mod_4626.get(0);
        mod_4627.put(0, t);
    endrule
    rule rule_5989;
        ChannelMessage t;
        t <- mod_4595.get(0);
        mod_4596.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4593.put(0, t);
        end
        if (i == 1) begin
            mod_4609.put(0, t);
        end
        if (i == 2) begin
            mod_4615.put(0, t);
        end
        if (i == 3) begin
            mod_4623.put(0, t);
        end
        if (i == 4) begin
            mod_4629.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_4597.get(0);
        end
        if (i == 3) begin
            t <- mod_4597.get(1);
        end
        if (i == 2) begin
            t <- mod_4597.get(2);
        end
        if (i == 1) begin
            t <- mod_4609.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6147 (Operation_IFC);
    Operation_IFC mod_4634_inner <- mkReshape(2, 64);
    Operation_IFC mod_4634 <- mkDebugOperation(mod_4634_inner, "mod_4634");
    Operation_IFC mod_4635_inner <- mkFlatten(1);
    Operation_IFC mod_4635 <- mkDebugOperation(mod_4635_inner, "mod_4635");
    Operation_IFC mod_4636_inner <- mkFlatten(2);
    Operation_IFC mod_4636 <- mkDebugOperation(mod_4636_inner, "mod_4636");
    Operation_IFC mod_4637_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4637 <- mkDebugOperation(mod_4637_inner, "mod_4637");
    Broadcast_IFC#(4) mod_4638_inner <- mkBroadcast(4);
    Operation_IFC mod_4638 <- mkDebugOperation(mod_4638_inner.op, "mod_4638");
    PMU_IFC mod_4639_bufferize <- mkPMU(2);
    Operation_IFC mod_4639_inner = mod_4639_bufferize.operation;
    Operation_IFC mod_4639 <- mkDebugOperation(mod_4639_inner, "mod_4639");
    Broadcast_IFC#(2) mod_4640_inner <- mkBroadcast(2);
    Operation_IFC mod_4640 <- mkDebugOperation(mod_4640_inner.op, "mod_4640");
    PMU_IFC mod_4641_bufferize <- mkPMU(1);
    Operation_IFC mod_4641_inner = mod_4641_bufferize.operation;
    Operation_IFC mod_4641 <- mkDebugOperation(mod_4641_inner, "mod_4641");
    Operation_IFC mod_4642_inner <- mkBinaryMap(1043, matmul_t_tile);
    Operation_IFC mod_4642 <- mkDebugOperation(mod_4642_inner, "mod_4642");
    Operation_IFC mod_4643_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4643 <- mkDebugOperation(mod_4643_inner, "mod_4643");
    Operation_IFC mod_4644_inner <- mkBinaryMap(1811, mul_tile);
    Operation_IFC mod_4644 <- mkDebugOperation(mod_4644_inner, "mod_4644");
    PMU_IFC mod_4645_bufferize <- mkPMU(1);
    Operation_IFC mod_4645_inner = mod_4645_bufferize.operation;
    Operation_IFC mod_4645 <- mkDebugOperation(mod_4645_inner, "mod_4645");
    Operation_IFC mod_4646_inner <- mkBinaryMap(2337, matmul_t_tile);
    Operation_IFC mod_4646 <- mkDebugOperation(mod_4646_inner, "mod_4646");
    Operation_IFC mod_4647_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4647 <- mkDebugOperation(mod_4647_inner, "mod_4647");
    Operation_IFC mod_4648_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4648 <- mkDebugOperation(mod_4648_inner, "mod_4648");
    Operation_IFC mod_4649_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4649 <- mkDebugOperation(mod_4649_inner, "mod_4649");
    Operation_IFC mod_4650_inner <- mkBinaryMap(2710, mul_tile);
    Operation_IFC mod_4650 <- mkDebugOperation(mod_4650_inner, "mod_4650");
    PMU_IFC mod_4651_bufferize <- mkPMU(1);
    Operation_IFC mod_4651_inner = mod_4651_bufferize.operation;
    Operation_IFC mod_4651 <- mkDebugOperation(mod_4651_inner, "mod_4651");
    PMU_IFC mod_4652_bufferize <- mkPMU(2);
    Operation_IFC mod_4652_inner = mod_4652_bufferize.operation;
    Operation_IFC mod_4652 <- mkDebugOperation(mod_4652_inner, "mod_4652");
    PMU_IFC mod_4653_bufferize <- mkPMU(2);
    Operation_IFC mod_4653_inner = mod_4653_bufferize.operation;
    Operation_IFC mod_4653 <- mkDebugOperation(mod_4653_inner, "mod_4653");
    Operation_IFC mod_4654_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4654 <- mkDebugOperation(mod_4654_inner, "mod_4654");
    Operation_IFC mod_4655_inner <- mkFlatten(1);
    Operation_IFC mod_4655 <- mkDebugOperation(mod_4655_inner, "mod_4655");
    Operation_IFC mod_4656_inner <- mkFlatten(0);
    Operation_IFC mod_4656 <- mkDebugOperation(mod_4656_inner, "mod_4656");
    Operation_IFC mod_4657_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4657 <- mkDebugOperation(mod_4657_inner, "mod_4657");
    Operation_IFC mod_4658_inner <- mkUnaryMap(1683, silu_tile);
    Operation_IFC mod_4658 <- mkDebugOperation(mod_4658_inner, "mod_4658");
    Operation_IFC mod_4659_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4659 <- mkDebugOperation(mod_4659_inner, "mod_4659");
    Operation_IFC mod_4660_inner <- mkBinaryMap(1555, matmul_t_tile);
    Operation_IFC mod_4660 <- mkDebugOperation(mod_4660_inner, "mod_4660");
    PMU_IFC mod_4661_bufferize <- mkPMU(2);
    Operation_IFC mod_4661_inner = mod_4661_bufferize.operation;
    Operation_IFC mod_4661 <- mkDebugOperation(mod_4661_inner, "mod_4661");
    Operation_IFC mod_4662_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4662 <- mkDebugOperation(mod_4662_inner, "mod_4662");
    Operation_IFC mod_4663_inner <- mkFlatten(1);
    Operation_IFC mod_4663 <- mkDebugOperation(mod_4663_inner, "mod_4663");
    Operation_IFC mod_4664_inner <- mkFlatten(0);
    Operation_IFC mod_4664 <- mkDebugOperation(mod_4664_inner, "mod_4664");
    PMU_IFC mod_4665_bufferize <- mkPMU(1);
    Operation_IFC mod_4665_inner = mod_4665_bufferize.operation;
    Operation_IFC mod_4665 <- mkDebugOperation(mod_4665_inner, "mod_4665");
    Operation_IFC mod_4666_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4666 <- mkDebugOperation(mod_4666_inner, "mod_4666");
    PMU_IFC mod_4667_bufferize <- mkPMU(2);
    Operation_IFC mod_4667_inner = mod_4667_bufferize.operation;
    Operation_IFC mod_4667 <- mkDebugOperation(mod_4667_inner, "mod_4667");
    Operation_IFC mod_4668_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4668 <- mkDebugOperation(mod_4668_inner, "mod_4668");
    Operation_IFC mod_4669_inner <- mkFlatten(1);
    Operation_IFC mod_4669 <- mkDebugOperation(mod_4669_inner, "mod_4669");
    Operation_IFC mod_4670_inner <- mkFlatten(0);
    Operation_IFC mod_4670 <- mkDebugOperation(mod_4670_inner, "mod_4670");
    Operation_IFC mod_4671_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4671 <- mkDebugOperation(mod_4671_inner, "mod_4671");
    Operation_IFC mod_4672_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4672 <- mkDebugOperation(mod_4672_inner, "mod_4672");
    PMU_IFC mod_4673_bufferize <- mkPMU(2);
    Operation_IFC mod_4673_inner = mod_4673_bufferize.operation;
    Operation_IFC mod_4673 <- mkDebugOperation(mod_4673_inner, "mod_4673");
    rule rule_5990;
        ChannelMessage t;
        t <- mod_4640.get(1);
        mod_4641.put(0, t);
    endrule
    rule rule_5991;
        ChannelMessage t;
        t <- mod_4637.get(0);
        mod_4673.put(0, t);
    endrule
    rule rule_5992;
        ChannelMessage t;
        t <- mod_4638.get(3);
        mod_4639.put(0, t);
    endrule
    rule rule_5993;
        ChannelMessage t;
        t <- mod_4651.get(1);
        mod_4649.put(1, t);
    endrule
    rule rule_5994;
        ChannelMessage t;
        t <- mod_4665.get(1);
        mod_4660.put(0, t);
    endrule
    rule rule_5995;
        ChannelMessage t;
        t <- mod_4645.get(0);
        mod_4657.put(0, t);
    endrule
    rule rule_5996;
        ChannelMessage t;
        t <- mod_4639.get(0);
        mod_4672.put(0, t);
    endrule
    rule rule_5997;
        ChannelMessage t;
        t <- mod_4673.get(0);
        mod_4673.put(1, t);
    endrule
    rule rule_5998;
        ChannelMessage t;
        t <- mod_4662.get(0);
        mod_4661.put(1, t);
    endrule
    rule rule_5999;
        ChannelMessage t;
        t <- mod_4653.get(0);
        mod_4654.put(0, t);
    endrule
    rule rule_6000;
        ChannelMessage t;
        t <- mod_4657.get(0);
        mod_4645.put(1, t);
    endrule
    rule rule_6001;
        ChannelMessage t;
        t <- mod_4663.get(0);
        mod_4661.put(0, t);
    endrule
    rule rule_6002;
        ChannelMessage t;
        t <- mod_4649.get(0);
        mod_4651.put(0, t);
    endrule
    rule rule_6003;
        ChannelMessage t;
        t <- mod_4671.get(0);
        mod_4641.put(1, t);
    endrule
    rule rule_6004;
        ChannelMessage t;
        t <- mod_4664.get(0);
        mod_4663.put(0, t);
    endrule
    rule rule_6005;
        ChannelMessage t;
        t <- mod_4670.get(0);
        mod_4669.put(0, t);
    endrule
    rule rule_6006;
        ChannelMessage t;
        t <- mod_4648.get(0);
        mod_4652.put(0, t);
    endrule
    rule rule_6007;
        ChannelMessage t;
        t <- mod_4644.get(0);
        mod_4645.put(0, t);
    endrule
    rule rule_6008;
        ChannelMessage t;
        t <- mod_4653.get(1);
        mod_4646.put(1, t);
    endrule
    rule rule_6009;
        ChannelMessage t;
        t <- mod_4660.get(0);
        mod_4659.put(0, t);
    endrule
    rule rule_6010;
        ChannelMessage t;
        t <- mod_4643.get(0);
        mod_4644.put(0, t);
    endrule
    rule rule_6011;
        ChannelMessage t;
        t <- mod_4635.get(0);
        mod_4636.put(0, t);
    endrule
    rule rule_6012;
        ChannelMessage t;
        t <- mod_4673.get(1);
        mod_4637.put(1, t);
    endrule
    rule rule_6013;
        ChannelMessage t;
        t <- mod_4647.get(0);
        mod_4648.put(0, t);
    endrule
    rule rule_6014;
        ChannelMessage t;
        t <- mod_4666.get(0);
        mod_4665.put(1, t);
    endrule
    rule rule_6015;
        ChannelMessage t;
        t <- mod_4651.get(0);
        mod_4651.put(1, t);
    endrule
    rule rule_6016;
        ChannelMessage t;
        t <- mod_4634.get(0);
        mod_4635.put(0, t);
    endrule
    rule rule_6017;
        ChannelMessage t;
        t <- mod_4652.get(1);
        mod_4648.put(1, t);
    endrule
    rule rule_6018;
        ChannelMessage t;
        t <- mod_4669.get(0);
        mod_4667.put(0, t);
    endrule
    rule rule_6019;
        ChannelMessage t;
        t <- mod_4658.get(0);
        mod_4644.put(1, t);
    endrule
    rule rule_6020;
        ChannelMessage t;
        t <- mod_4665.get(0);
        mod_4666.put(0, t);
    endrule
    rule rule_6021;
        ChannelMessage t;
        t <- mod_4667.get(1);
        mod_4642.put(1, t);
    endrule
    rule rule_6022;
        ChannelMessage t;
        t <- mod_4640.get(0);
        mod_4665.put(0, t);
    endrule
    rule rule_6023;
        ChannelMessage t;
        t <- mod_4668.get(0);
        mod_4667.put(1, t);
    endrule
    rule rule_6024;
        ChannelMessage t;
        t <- mod_4655.get(0);
        mod_4653.put(0, t);
    endrule
    rule rule_6025;
        ChannelMessage t;
        t <- mod_4646.get(0);
        mod_4647.put(0, t);
    endrule
    rule rule_6026;
        ChannelMessage t;
        t <- mod_4637.get(1);
        mod_4638.put(0, t);
    endrule
    rule rule_6027;
        ChannelMessage t;
        t <- mod_4636.get(0);
        mod_4637.put(0, t);
    endrule
    rule rule_6028;
        ChannelMessage t;
        t <- mod_4652.get(0);
        mod_4652.put(1, t);
    endrule
    rule rule_6029;
        ChannelMessage t;
        t <- mod_4661.get(1);
        mod_4660.put(1, t);
    endrule
    rule rule_6030;
        ChannelMessage t;
        t <- mod_4661.get(0);
        mod_4662.put(0, t);
    endrule
    rule rule_6031;
        ChannelMessage t;
        t <- mod_4642.get(0);
        mod_4643.put(0, t);
    endrule
    rule rule_6032;
        ChannelMessage t;
        t <- mod_4645.get(1);
        mod_4646.put(0, t);
    endrule
    rule rule_6033;
        ChannelMessage t;
        t <- mod_4654.get(0);
        mod_4653.put(1, t);
    endrule
    rule rule_6034;
        ChannelMessage t;
        t <- mod_4667.get(0);
        mod_4668.put(0, t);
    endrule
    rule rule_6035;
        ChannelMessage t;
        t <- mod_4656.get(0);
        mod_4655.put(0, t);
    endrule
    rule rule_6036;
        ChannelMessage t;
        t <- mod_4672.get(0);
        mod_4639.put(1, t);
    endrule
    rule rule_6037;
        ChannelMessage t;
        t <- mod_4659.get(0);
        mod_4658.put(0, t);
    endrule
    rule rule_6038;
        ChannelMessage t;
        t <- mod_4648.get(1);
        mod_4649.put(0, t);
    endrule
    rule rule_6039;
        ChannelMessage t;
        t <- mod_4641.get(1);
        mod_4642.put(0, t);
    endrule
    rule rule_6040;
        ChannelMessage t;
        t <- mod_4639.get(1);
        mod_4640.put(0, t);
    endrule
    rule rule_6041;
        ChannelMessage t;
        t <- mod_4649.get(1);
        mod_4650.put(1, t);
    endrule
    rule rule_6042;
        ChannelMessage t;
        t <- mod_4641.get(0);
        mod_4671.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4634.put(0, t);
        end
        if (i == 1) begin
            mod_4650.put(0, t);
        end
        if (i == 2) begin
            mod_4656.put(0, t);
        end
        if (i == 3) begin
            mod_4664.put(0, t);
        end
        if (i == 4) begin
            mod_4670.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_4638.get(0);
        end
        if (i == 3) begin
            t <- mod_4638.get(1);
        end
        if (i == 2) begin
            t <- mod_4638.get(2);
        end
        if (i == 0) begin
            t <- mod_4650.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6148 (Operation_IFC);
    Operation_IFC mod_4675_inner <- mkReshape(2, 64);
    Operation_IFC mod_4675 <- mkDebugOperation(mod_4675_inner, "mod_4675");
    Operation_IFC mod_4676_inner <- mkFlatten(1);
    Operation_IFC mod_4676 <- mkDebugOperation(mod_4676_inner, "mod_4676");
    Operation_IFC mod_4677_inner <- mkFlatten(2);
    Operation_IFC mod_4677 <- mkDebugOperation(mod_4677_inner, "mod_4677");
    Operation_IFC mod_4678_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4678 <- mkDebugOperation(mod_4678_inner, "mod_4678");
    Broadcast_IFC#(4) mod_4679_inner <- mkBroadcast(4);
    Operation_IFC mod_4679 <- mkDebugOperation(mod_4679_inner.op, "mod_4679");
    PMU_IFC mod_4680_bufferize <- mkPMU(2);
    Operation_IFC mod_4680_inner = mod_4680_bufferize.operation;
    Operation_IFC mod_4680 <- mkDebugOperation(mod_4680_inner, "mod_4680");
    Broadcast_IFC#(2) mod_4681_inner <- mkBroadcast(2);
    Operation_IFC mod_4681 <- mkDebugOperation(mod_4681_inner.op, "mod_4681");
    PMU_IFC mod_4682_bufferize <- mkPMU(1);
    Operation_IFC mod_4682_inner = mod_4682_bufferize.operation;
    Operation_IFC mod_4682 <- mkDebugOperation(mod_4682_inner, "mod_4682");
    Operation_IFC mod_4683_inner <- mkBinaryMap(1042, matmul_t_tile);
    Operation_IFC mod_4683 <- mkDebugOperation(mod_4683_inner, "mod_4683");
    Operation_IFC mod_4684_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4684 <- mkDebugOperation(mod_4684_inner, "mod_4684");
    Operation_IFC mod_4685_inner <- mkBinaryMap(1810, mul_tile);
    Operation_IFC mod_4685 <- mkDebugOperation(mod_4685_inner, "mod_4685");
    PMU_IFC mod_4686_bufferize <- mkPMU(1);
    Operation_IFC mod_4686_inner = mod_4686_bufferize.operation;
    Operation_IFC mod_4686 <- mkDebugOperation(mod_4686_inner, "mod_4686");
    Operation_IFC mod_4687_inner <- mkBinaryMap(2335, matmul_t_tile);
    Operation_IFC mod_4687 <- mkDebugOperation(mod_4687_inner, "mod_4687");
    Operation_IFC mod_4688_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4688 <- mkDebugOperation(mod_4688_inner, "mod_4688");
    Operation_IFC mod_4689_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4689 <- mkDebugOperation(mod_4689_inner, "mod_4689");
    Operation_IFC mod_4690_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4690 <- mkDebugOperation(mod_4690_inner, "mod_4690");
    Operation_IFC mod_4691_inner <- mkBinaryMap(2709, mul_tile);
    Operation_IFC mod_4691 <- mkDebugOperation(mod_4691_inner, "mod_4691");
    PMU_IFC mod_4692_bufferize <- mkPMU(1);
    Operation_IFC mod_4692_inner = mod_4692_bufferize.operation;
    Operation_IFC mod_4692 <- mkDebugOperation(mod_4692_inner, "mod_4692");
    PMU_IFC mod_4693_bufferize <- mkPMU(2);
    Operation_IFC mod_4693_inner = mod_4693_bufferize.operation;
    Operation_IFC mod_4693 <- mkDebugOperation(mod_4693_inner, "mod_4693");
    PMU_IFC mod_4694_bufferize <- mkPMU(2);
    Operation_IFC mod_4694_inner = mod_4694_bufferize.operation;
    Operation_IFC mod_4694 <- mkDebugOperation(mod_4694_inner, "mod_4694");
    Operation_IFC mod_4695_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4695 <- mkDebugOperation(mod_4695_inner, "mod_4695");
    Operation_IFC mod_4696_inner <- mkFlatten(1);
    Operation_IFC mod_4696 <- mkDebugOperation(mod_4696_inner, "mod_4696");
    Operation_IFC mod_4697_inner <- mkFlatten(0);
    Operation_IFC mod_4697 <- mkDebugOperation(mod_4697_inner, "mod_4697");
    Operation_IFC mod_4698_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4698 <- mkDebugOperation(mod_4698_inner, "mod_4698");
    Operation_IFC mod_4699_inner <- mkUnaryMap(1682, silu_tile);
    Operation_IFC mod_4699 <- mkDebugOperation(mod_4699_inner, "mod_4699");
    Operation_IFC mod_4700_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4700 <- mkDebugOperation(mod_4700_inner, "mod_4700");
    Operation_IFC mod_4701_inner <- mkBinaryMap(1554, matmul_t_tile);
    Operation_IFC mod_4701 <- mkDebugOperation(mod_4701_inner, "mod_4701");
    PMU_IFC mod_4702_bufferize <- mkPMU(2);
    Operation_IFC mod_4702_inner = mod_4702_bufferize.operation;
    Operation_IFC mod_4702 <- mkDebugOperation(mod_4702_inner, "mod_4702");
    Operation_IFC mod_4703_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4703 <- mkDebugOperation(mod_4703_inner, "mod_4703");
    Operation_IFC mod_4704_inner <- mkFlatten(1);
    Operation_IFC mod_4704 <- mkDebugOperation(mod_4704_inner, "mod_4704");
    Operation_IFC mod_4705_inner <- mkFlatten(0);
    Operation_IFC mod_4705 <- mkDebugOperation(mod_4705_inner, "mod_4705");
    PMU_IFC mod_4706_bufferize <- mkPMU(1);
    Operation_IFC mod_4706_inner = mod_4706_bufferize.operation;
    Operation_IFC mod_4706 <- mkDebugOperation(mod_4706_inner, "mod_4706");
    Operation_IFC mod_4707_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4707 <- mkDebugOperation(mod_4707_inner, "mod_4707");
    PMU_IFC mod_4708_bufferize <- mkPMU(2);
    Operation_IFC mod_4708_inner = mod_4708_bufferize.operation;
    Operation_IFC mod_4708 <- mkDebugOperation(mod_4708_inner, "mod_4708");
    Operation_IFC mod_4709_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4709 <- mkDebugOperation(mod_4709_inner, "mod_4709");
    Operation_IFC mod_4710_inner <- mkFlatten(1);
    Operation_IFC mod_4710 <- mkDebugOperation(mod_4710_inner, "mod_4710");
    Operation_IFC mod_4711_inner <- mkFlatten(0);
    Operation_IFC mod_4711 <- mkDebugOperation(mod_4711_inner, "mod_4711");
    Operation_IFC mod_4712_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4712 <- mkDebugOperation(mod_4712_inner, "mod_4712");
    Operation_IFC mod_4713_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4713 <- mkDebugOperation(mod_4713_inner, "mod_4713");
    PMU_IFC mod_4714_bufferize <- mkPMU(2);
    Operation_IFC mod_4714_inner = mod_4714_bufferize.operation;
    Operation_IFC mod_4714 <- mkDebugOperation(mod_4714_inner, "mod_4714");
    rule rule_6043;
        ChannelMessage t;
        t <- mod_4706.get(1);
        mod_4701.put(0, t);
    endrule
    rule rule_6044;
        ChannelMessage t;
        t <- mod_4684.get(0);
        mod_4685.put(0, t);
    endrule
    rule rule_6045;
        ChannelMessage t;
        t <- mod_4676.get(0);
        mod_4677.put(0, t);
    endrule
    rule rule_6046;
        ChannelMessage t;
        t <- mod_4682.get(0);
        mod_4712.put(0, t);
    endrule
    rule rule_6047;
        ChannelMessage t;
        t <- mod_4687.get(0);
        mod_4688.put(0, t);
    endrule
    rule rule_6048;
        ChannelMessage t;
        t <- mod_4708.get(0);
        mod_4709.put(0, t);
    endrule
    rule rule_6049;
        ChannelMessage t;
        t <- mod_4681.get(1);
        mod_4682.put(0, t);
    endrule
    rule rule_6050;
        ChannelMessage t;
        t <- mod_4696.get(0);
        mod_4694.put(0, t);
    endrule
    rule rule_6051;
        ChannelMessage t;
        t <- mod_4689.get(1);
        mod_4690.put(0, t);
    endrule
    rule rule_6052;
        ChannelMessage t;
        t <- mod_4693.get(0);
        mod_4693.put(1, t);
    endrule
    rule rule_6053;
        ChannelMessage t;
        t <- mod_4694.get(0);
        mod_4695.put(0, t);
    endrule
    rule rule_6054;
        ChannelMessage t;
        t <- mod_4692.get(0);
        mod_4692.put(1, t);
    endrule
    rule rule_6055;
        ChannelMessage t;
        t <- mod_4688.get(0);
        mod_4689.put(0, t);
    endrule
    rule rule_6056;
        ChannelMessage t;
        t <- mod_4703.get(0);
        mod_4702.put(1, t);
    endrule
    rule rule_6057;
        ChannelMessage t;
        t <- mod_4705.get(0);
        mod_4704.put(0, t);
    endrule
    rule rule_6058;
        ChannelMessage t;
        t <- mod_4706.get(0);
        mod_4707.put(0, t);
    endrule
    rule rule_6059;
        ChannelMessage t;
        t <- mod_4690.get(0);
        mod_4692.put(0, t);
    endrule
    rule rule_6060;
        ChannelMessage t;
        t <- mod_4700.get(0);
        mod_4699.put(0, t);
    endrule
    rule rule_6061;
        ChannelMessage t;
        t <- mod_4677.get(0);
        mod_4678.put(0, t);
    endrule
    rule rule_6062;
        ChannelMessage t;
        t <- mod_4682.get(1);
        mod_4683.put(0, t);
    endrule
    rule rule_6063;
        ChannelMessage t;
        t <- mod_4710.get(0);
        mod_4708.put(0, t);
    endrule
    rule rule_6064;
        ChannelMessage t;
        t <- mod_4686.get(0);
        mod_4698.put(0, t);
    endrule
    rule rule_6065;
        ChannelMessage t;
        t <- mod_4679.get(3);
        mod_4680.put(0, t);
    endrule
    rule rule_6066;
        ChannelMessage t;
        t <- mod_4680.get(0);
        mod_4713.put(0, t);
    endrule
    rule rule_6067;
        ChannelMessage t;
        t <- mod_4707.get(0);
        mod_4706.put(1, t);
    endrule
    rule rule_6068;
        ChannelMessage t;
        t <- mod_4708.get(1);
        mod_4683.put(1, t);
    endrule
    rule rule_6069;
        ChannelMessage t;
        t <- mod_4713.get(0);
        mod_4680.put(1, t);
    endrule
    rule rule_6070;
        ChannelMessage t;
        t <- mod_4693.get(1);
        mod_4689.put(1, t);
    endrule
    rule rule_6071;
        ChannelMessage t;
        t <- mod_4692.get(1);
        mod_4690.put(1, t);
    endrule
    rule rule_6072;
        ChannelMessage t;
        t <- mod_4683.get(0);
        mod_4684.put(0, t);
    endrule
    rule rule_6073;
        ChannelMessage t;
        t <- mod_4702.get(1);
        mod_4701.put(1, t);
    endrule
    rule rule_6074;
        ChannelMessage t;
        t <- mod_4678.get(0);
        mod_4714.put(0, t);
    endrule
    rule rule_6075;
        ChannelMessage t;
        t <- mod_4709.get(0);
        mod_4708.put(1, t);
    endrule
    rule rule_6076;
        ChannelMessage t;
        t <- mod_4695.get(0);
        mod_4694.put(1, t);
    endrule
    rule rule_6077;
        ChannelMessage t;
        t <- mod_4678.get(1);
        mod_4679.put(0, t);
    endrule
    rule rule_6078;
        ChannelMessage t;
        t <- mod_4689.get(0);
        mod_4693.put(0, t);
    endrule
    rule rule_6079;
        ChannelMessage t;
        t <- mod_4699.get(0);
        mod_4685.put(1, t);
    endrule
    rule rule_6080;
        ChannelMessage t;
        t <- mod_4701.get(0);
        mod_4700.put(0, t);
    endrule
    rule rule_6081;
        ChannelMessage t;
        t <- mod_4697.get(0);
        mod_4696.put(0, t);
    endrule
    rule rule_6082;
        ChannelMessage t;
        t <- mod_4712.get(0);
        mod_4682.put(1, t);
    endrule
    rule rule_6083;
        ChannelMessage t;
        t <- mod_4685.get(0);
        mod_4686.put(0, t);
    endrule
    rule rule_6084;
        ChannelMessage t;
        t <- mod_4711.get(0);
        mod_4710.put(0, t);
    endrule
    rule rule_6085;
        ChannelMessage t;
        t <- mod_4680.get(1);
        mod_4681.put(0, t);
    endrule
    rule rule_6086;
        ChannelMessage t;
        t <- mod_4704.get(0);
        mod_4702.put(0, t);
    endrule
    rule rule_6087;
        ChannelMessage t;
        t <- mod_4690.get(1);
        mod_4691.put(1, t);
    endrule
    rule rule_6088;
        ChannelMessage t;
        t <- mod_4714.get(1);
        mod_4678.put(1, t);
    endrule
    rule rule_6089;
        ChannelMessage t;
        t <- mod_4675.get(0);
        mod_4676.put(0, t);
    endrule
    rule rule_6090;
        ChannelMessage t;
        t <- mod_4714.get(0);
        mod_4714.put(1, t);
    endrule
    rule rule_6091;
        ChannelMessage t;
        t <- mod_4694.get(1);
        mod_4687.put(1, t);
    endrule
    rule rule_6092;
        ChannelMessage t;
        t <- mod_4698.get(0);
        mod_4686.put(1, t);
    endrule
    rule rule_6093;
        ChannelMessage t;
        t <- mod_4681.get(0);
        mod_4706.put(0, t);
    endrule
    rule rule_6094;
        ChannelMessage t;
        t <- mod_4686.get(1);
        mod_4687.put(0, t);
    endrule
    rule rule_6095;
        ChannelMessage t;
        t <- mod_4702.get(0);
        mod_4703.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4675.put(0, t);
        end
        if (i == 1) begin
            mod_4691.put(0, t);
        end
        if (i == 2) begin
            mod_4697.put(0, t);
        end
        if (i == 3) begin
            mod_4705.put(0, t);
        end
        if (i == 4) begin
            mod_4711.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_4679.get(0);
        end
        if (i == 1) begin
            t <- mod_4679.get(1);
        end
        if (i == 3) begin
            t <- mod_4679.get(2);
        end
        if (i == 2) begin
            t <- mod_4691.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6149 (Operation_IFC);
    Operation_IFC mod_4716_inner <- mkReshape(2, 64);
    Operation_IFC mod_4716 <- mkDebugOperation(mod_4716_inner, "mod_4716");
    Operation_IFC mod_4717_inner <- mkFlatten(1);
    Operation_IFC mod_4717 <- mkDebugOperation(mod_4717_inner, "mod_4717");
    Operation_IFC mod_4718_inner <- mkFlatten(2);
    Operation_IFC mod_4718 <- mkDebugOperation(mod_4718_inner, "mod_4718");
    Operation_IFC mod_4719_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4719 <- mkDebugOperation(mod_4719_inner, "mod_4719");
    Broadcast_IFC#(4) mod_4720_inner <- mkBroadcast(4);
    Operation_IFC mod_4720 <- mkDebugOperation(mod_4720_inner.op, "mod_4720");
    PMU_IFC mod_4721_bufferize <- mkPMU(2);
    Operation_IFC mod_4721_inner = mod_4721_bufferize.operation;
    Operation_IFC mod_4721 <- mkDebugOperation(mod_4721_inner, "mod_4721");
    Broadcast_IFC#(2) mod_4722_inner <- mkBroadcast(2);
    Operation_IFC mod_4722 <- mkDebugOperation(mod_4722_inner.op, "mod_4722");
    PMU_IFC mod_4723_bufferize <- mkPMU(1);
    Operation_IFC mod_4723_inner = mod_4723_bufferize.operation;
    Operation_IFC mod_4723 <- mkDebugOperation(mod_4723_inner, "mod_4723");
    Operation_IFC mod_4724_inner <- mkBinaryMap(1041, matmul_t_tile);
    Operation_IFC mod_4724 <- mkDebugOperation(mod_4724_inner, "mod_4724");
    Operation_IFC mod_4725_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4725 <- mkDebugOperation(mod_4725_inner, "mod_4725");
    Operation_IFC mod_4726_inner <- mkBinaryMap(1809, mul_tile);
    Operation_IFC mod_4726 <- mkDebugOperation(mod_4726_inner, "mod_4726");
    PMU_IFC mod_4727_bufferize <- mkPMU(1);
    Operation_IFC mod_4727_inner = mod_4727_bufferize.operation;
    Operation_IFC mod_4727 <- mkDebugOperation(mod_4727_inner, "mod_4727");
    Operation_IFC mod_4728_inner <- mkBinaryMap(2333, matmul_t_tile);
    Operation_IFC mod_4728 <- mkDebugOperation(mod_4728_inner, "mod_4728");
    Operation_IFC mod_4729_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4729 <- mkDebugOperation(mod_4729_inner, "mod_4729");
    Operation_IFC mod_4730_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4730 <- mkDebugOperation(mod_4730_inner, "mod_4730");
    Operation_IFC mod_4731_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4731 <- mkDebugOperation(mod_4731_inner, "mod_4731");
    Operation_IFC mod_4732_inner <- mkBinaryMap(2708, mul_tile);
    Operation_IFC mod_4732 <- mkDebugOperation(mod_4732_inner, "mod_4732");
    PMU_IFC mod_4733_bufferize <- mkPMU(1);
    Operation_IFC mod_4733_inner = mod_4733_bufferize.operation;
    Operation_IFC mod_4733 <- mkDebugOperation(mod_4733_inner, "mod_4733");
    PMU_IFC mod_4734_bufferize <- mkPMU(2);
    Operation_IFC mod_4734_inner = mod_4734_bufferize.operation;
    Operation_IFC mod_4734 <- mkDebugOperation(mod_4734_inner, "mod_4734");
    PMU_IFC mod_4735_bufferize <- mkPMU(2);
    Operation_IFC mod_4735_inner = mod_4735_bufferize.operation;
    Operation_IFC mod_4735 <- mkDebugOperation(mod_4735_inner, "mod_4735");
    Operation_IFC mod_4736_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4736 <- mkDebugOperation(mod_4736_inner, "mod_4736");
    Operation_IFC mod_4737_inner <- mkFlatten(1);
    Operation_IFC mod_4737 <- mkDebugOperation(mod_4737_inner, "mod_4737");
    Operation_IFC mod_4738_inner <- mkFlatten(0);
    Operation_IFC mod_4738 <- mkDebugOperation(mod_4738_inner, "mod_4738");
    Operation_IFC mod_4739_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4739 <- mkDebugOperation(mod_4739_inner, "mod_4739");
    Operation_IFC mod_4740_inner <- mkUnaryMap(1681, silu_tile);
    Operation_IFC mod_4740 <- mkDebugOperation(mod_4740_inner, "mod_4740");
    Operation_IFC mod_4741_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4741 <- mkDebugOperation(mod_4741_inner, "mod_4741");
    Operation_IFC mod_4742_inner <- mkBinaryMap(1553, matmul_t_tile);
    Operation_IFC mod_4742 <- mkDebugOperation(mod_4742_inner, "mod_4742");
    PMU_IFC mod_4743_bufferize <- mkPMU(2);
    Operation_IFC mod_4743_inner = mod_4743_bufferize.operation;
    Operation_IFC mod_4743 <- mkDebugOperation(mod_4743_inner, "mod_4743");
    Operation_IFC mod_4744_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4744 <- mkDebugOperation(mod_4744_inner, "mod_4744");
    Operation_IFC mod_4745_inner <- mkFlatten(1);
    Operation_IFC mod_4745 <- mkDebugOperation(mod_4745_inner, "mod_4745");
    Operation_IFC mod_4746_inner <- mkFlatten(0);
    Operation_IFC mod_4746 <- mkDebugOperation(mod_4746_inner, "mod_4746");
    PMU_IFC mod_4747_bufferize <- mkPMU(1);
    Operation_IFC mod_4747_inner = mod_4747_bufferize.operation;
    Operation_IFC mod_4747 <- mkDebugOperation(mod_4747_inner, "mod_4747");
    Operation_IFC mod_4748_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4748 <- mkDebugOperation(mod_4748_inner, "mod_4748");
    PMU_IFC mod_4749_bufferize <- mkPMU(2);
    Operation_IFC mod_4749_inner = mod_4749_bufferize.operation;
    Operation_IFC mod_4749 <- mkDebugOperation(mod_4749_inner, "mod_4749");
    Operation_IFC mod_4750_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4750 <- mkDebugOperation(mod_4750_inner, "mod_4750");
    Operation_IFC mod_4751_inner <- mkFlatten(1);
    Operation_IFC mod_4751 <- mkDebugOperation(mod_4751_inner, "mod_4751");
    Operation_IFC mod_4752_inner <- mkFlatten(0);
    Operation_IFC mod_4752 <- mkDebugOperation(mod_4752_inner, "mod_4752");
    Operation_IFC mod_4753_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4753 <- mkDebugOperation(mod_4753_inner, "mod_4753");
    Operation_IFC mod_4754_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4754 <- mkDebugOperation(mod_4754_inner, "mod_4754");
    PMU_IFC mod_4755_bufferize <- mkPMU(2);
    Operation_IFC mod_4755_inner = mod_4755_bufferize.operation;
    Operation_IFC mod_4755 <- mkDebugOperation(mod_4755_inner, "mod_4755");
    rule rule_6096;
        ChannelMessage t;
        t <- mod_4755.get(0);
        mod_4755.put(1, t);
    endrule
    rule rule_6097;
        ChannelMessage t;
        t <- mod_4728.get(0);
        mod_4729.put(0, t);
    endrule
    rule rule_6098;
        ChannelMessage t;
        t <- mod_4738.get(0);
        mod_4737.put(0, t);
    endrule
    rule rule_6099;
        ChannelMessage t;
        t <- mod_4750.get(0);
        mod_4749.put(1, t);
    endrule
    rule rule_6100;
        ChannelMessage t;
        t <- mod_4727.get(0);
        mod_4739.put(0, t);
    endrule
    rule rule_6101;
        ChannelMessage t;
        t <- mod_4743.get(0);
        mod_4744.put(0, t);
    endrule
    rule rule_6102;
        ChannelMessage t;
        t <- mod_4730.get(1);
        mod_4731.put(0, t);
    endrule
    rule rule_6103;
        ChannelMessage t;
        t <- mod_4740.get(0);
        mod_4726.put(1, t);
    endrule
    rule rule_6104;
        ChannelMessage t;
        t <- mod_4735.get(1);
        mod_4728.put(1, t);
    endrule
    rule rule_6105;
        ChannelMessage t;
        t <- mod_4749.get(1);
        mod_4724.put(1, t);
    endrule
    rule rule_6106;
        ChannelMessage t;
        t <- mod_4722.get(1);
        mod_4723.put(0, t);
    endrule
    rule rule_6107;
        ChannelMessage t;
        t <- mod_4747.get(0);
        mod_4748.put(0, t);
    endrule
    rule rule_6108;
        ChannelMessage t;
        t <- mod_4731.get(0);
        mod_4733.put(0, t);
    endrule
    rule rule_6109;
        ChannelMessage t;
        t <- mod_4745.get(0);
        mod_4743.put(0, t);
    endrule
    rule rule_6110;
        ChannelMessage t;
        t <- mod_4755.get(1);
        mod_4719.put(1, t);
    endrule
    rule rule_6111;
        ChannelMessage t;
        t <- mod_4747.get(1);
        mod_4742.put(0, t);
    endrule
    rule rule_6112;
        ChannelMessage t;
        t <- mod_4748.get(0);
        mod_4747.put(1, t);
    endrule
    rule rule_6113;
        ChannelMessage t;
        t <- mod_4719.get(0);
        mod_4755.put(0, t);
    endrule
    rule rule_6114;
        ChannelMessage t;
        t <- mod_4719.get(1);
        mod_4720.put(0, t);
    endrule
    rule rule_6115;
        ChannelMessage t;
        t <- mod_4741.get(0);
        mod_4740.put(0, t);
    endrule
    rule rule_6116;
        ChannelMessage t;
        t <- mod_4730.get(0);
        mod_4734.put(0, t);
    endrule
    rule rule_6117;
        ChannelMessage t;
        t <- mod_4746.get(0);
        mod_4745.put(0, t);
    endrule
    rule rule_6118;
        ChannelMessage t;
        t <- mod_4752.get(0);
        mod_4751.put(0, t);
    endrule
    rule rule_6119;
        ChannelMessage t;
        t <- mod_4736.get(0);
        mod_4735.put(1, t);
    endrule
    rule rule_6120;
        ChannelMessage t;
        t <- mod_4723.get(1);
        mod_4724.put(0, t);
    endrule
    rule rule_6121;
        ChannelMessage t;
        t <- mod_4733.get(0);
        mod_4733.put(1, t);
    endrule
    rule rule_6122;
        ChannelMessage t;
        t <- mod_4722.get(0);
        mod_4747.put(0, t);
    endrule
    rule rule_6123;
        ChannelMessage t;
        t <- mod_4734.get(0);
        mod_4734.put(1, t);
    endrule
    rule rule_6124;
        ChannelMessage t;
        t <- mod_4753.get(0);
        mod_4723.put(1, t);
    endrule
    rule rule_6125;
        ChannelMessage t;
        t <- mod_4743.get(1);
        mod_4742.put(1, t);
    endrule
    rule rule_6126;
        ChannelMessage t;
        t <- mod_4720.get(3);
        mod_4721.put(0, t);
    endrule
    rule rule_6127;
        ChannelMessage t;
        t <- mod_4725.get(0);
        mod_4726.put(0, t);
    endrule
    rule rule_6128;
        ChannelMessage t;
        t <- mod_4723.get(0);
        mod_4753.put(0, t);
    endrule
    rule rule_6129;
        ChannelMessage t;
        t <- mod_4721.get(0);
        mod_4754.put(0, t);
    endrule
    rule rule_6130;
        ChannelMessage t;
        t <- mod_4727.get(1);
        mod_4728.put(0, t);
    endrule
    rule rule_6131;
        ChannelMessage t;
        t <- mod_4744.get(0);
        mod_4743.put(1, t);
    endrule
    rule rule_6132;
        ChannelMessage t;
        t <- mod_4718.get(0);
        mod_4719.put(0, t);
    endrule
    rule rule_6133;
        ChannelMessage t;
        t <- mod_4754.get(0);
        mod_4721.put(1, t);
    endrule
    rule rule_6134;
        ChannelMessage t;
        t <- mod_4737.get(0);
        mod_4735.put(0, t);
    endrule
    rule rule_6135;
        ChannelMessage t;
        t <- mod_4721.get(1);
        mod_4722.put(0, t);
    endrule
    rule rule_6136;
        ChannelMessage t;
        t <- mod_4733.get(1);
        mod_4731.put(1, t);
    endrule
    rule rule_6137;
        ChannelMessage t;
        t <- mod_4751.get(0);
        mod_4749.put(0, t);
    endrule
    rule rule_6138;
        ChannelMessage t;
        t <- mod_4735.get(0);
        mod_4736.put(0, t);
    endrule
    rule rule_6139;
        ChannelMessage t;
        t <- mod_4724.get(0);
        mod_4725.put(0, t);
    endrule
    rule rule_6140;
        ChannelMessage t;
        t <- mod_4731.get(1);
        mod_4732.put(1, t);
    endrule
    rule rule_6141;
        ChannelMessage t;
        t <- mod_4749.get(0);
        mod_4750.put(0, t);
    endrule
    rule rule_6142;
        ChannelMessage t;
        t <- mod_4729.get(0);
        mod_4730.put(0, t);
    endrule
    rule rule_6143;
        ChannelMessage t;
        t <- mod_4717.get(0);
        mod_4718.put(0, t);
    endrule
    rule rule_6144;
        ChannelMessage t;
        t <- mod_4726.get(0);
        mod_4727.put(0, t);
    endrule
    rule rule_6145;
        ChannelMessage t;
        t <- mod_4716.get(0);
        mod_4717.put(0, t);
    endrule
    rule rule_6146;
        ChannelMessage t;
        t <- mod_4734.get(1);
        mod_4730.put(1, t);
    endrule
    rule rule_6147;
        ChannelMessage t;
        t <- mod_4742.get(0);
        mod_4741.put(0, t);
    endrule
    rule rule_6148;
        ChannelMessage t;
        t <- mod_4739.get(0);
        mod_4727.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4716.put(0, t);
        end
        if (i == 1) begin
            mod_4732.put(0, t);
        end
        if (i == 2) begin
            mod_4738.put(0, t);
        end
        if (i == 3) begin
            mod_4746.put(0, t);
        end
        if (i == 4) begin
            mod_4752.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_4720.get(0);
        end
        if (i == 2) begin
            t <- mod_4720.get(1);
        end
        if (i == 1) begin
            t <- mod_4720.get(2);
        end
        if (i == 3) begin
            t <- mod_4732.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6150 (Operation_IFC);
    Operation_IFC mod_4757_inner <- mkReshape(2, 64);
    Operation_IFC mod_4757 <- mkDebugOperation(mod_4757_inner, "mod_4757");
    Operation_IFC mod_4758_inner <- mkFlatten(1);
    Operation_IFC mod_4758 <- mkDebugOperation(mod_4758_inner, "mod_4758");
    Operation_IFC mod_4759_inner <- mkFlatten(2);
    Operation_IFC mod_4759 <- mkDebugOperation(mod_4759_inner, "mod_4759");
    Operation_IFC mod_4760_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4760 <- mkDebugOperation(mod_4760_inner, "mod_4760");
    Broadcast_IFC#(4) mod_4761_inner <- mkBroadcast(4);
    Operation_IFC mod_4761 <- mkDebugOperation(mod_4761_inner.op, "mod_4761");
    PMU_IFC mod_4762_bufferize <- mkPMU(2);
    Operation_IFC mod_4762_inner = mod_4762_bufferize.operation;
    Operation_IFC mod_4762 <- mkDebugOperation(mod_4762_inner, "mod_4762");
    Broadcast_IFC#(2) mod_4763_inner <- mkBroadcast(2);
    Operation_IFC mod_4763 <- mkDebugOperation(mod_4763_inner.op, "mod_4763");
    PMU_IFC mod_4764_bufferize <- mkPMU(1);
    Operation_IFC mod_4764_inner = mod_4764_bufferize.operation;
    Operation_IFC mod_4764 <- mkDebugOperation(mod_4764_inner, "mod_4764");
    Operation_IFC mod_4765_inner <- mkBinaryMap(1040, matmul_t_tile);
    Operation_IFC mod_4765 <- mkDebugOperation(mod_4765_inner, "mod_4765");
    Operation_IFC mod_4766_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4766 <- mkDebugOperation(mod_4766_inner, "mod_4766");
    Operation_IFC mod_4767_inner <- mkBinaryMap(1808, mul_tile);
    Operation_IFC mod_4767 <- mkDebugOperation(mod_4767_inner, "mod_4767");
    PMU_IFC mod_4768_bufferize <- mkPMU(1);
    Operation_IFC mod_4768_inner = mod_4768_bufferize.operation;
    Operation_IFC mod_4768 <- mkDebugOperation(mod_4768_inner, "mod_4768");
    Operation_IFC mod_4769_inner <- mkBinaryMap(2331, matmul_t_tile);
    Operation_IFC mod_4769 <- mkDebugOperation(mod_4769_inner, "mod_4769");
    Operation_IFC mod_4770_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4770 <- mkDebugOperation(mod_4770_inner, "mod_4770");
    Operation_IFC mod_4771_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4771 <- mkDebugOperation(mod_4771_inner, "mod_4771");
    Operation_IFC mod_4772_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4772 <- mkDebugOperation(mod_4772_inner, "mod_4772");
    Operation_IFC mod_4773_inner <- mkBinaryMap(2707, mul_tile);
    Operation_IFC mod_4773 <- mkDebugOperation(mod_4773_inner, "mod_4773");
    PMU_IFC mod_4774_bufferize <- mkPMU(1);
    Operation_IFC mod_4774_inner = mod_4774_bufferize.operation;
    Operation_IFC mod_4774 <- mkDebugOperation(mod_4774_inner, "mod_4774");
    PMU_IFC mod_4775_bufferize <- mkPMU(2);
    Operation_IFC mod_4775_inner = mod_4775_bufferize.operation;
    Operation_IFC mod_4775 <- mkDebugOperation(mod_4775_inner, "mod_4775");
    PMU_IFC mod_4776_bufferize <- mkPMU(2);
    Operation_IFC mod_4776_inner = mod_4776_bufferize.operation;
    Operation_IFC mod_4776 <- mkDebugOperation(mod_4776_inner, "mod_4776");
    Operation_IFC mod_4777_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4777 <- mkDebugOperation(mod_4777_inner, "mod_4777");
    Operation_IFC mod_4778_inner <- mkFlatten(1);
    Operation_IFC mod_4778 <- mkDebugOperation(mod_4778_inner, "mod_4778");
    Operation_IFC mod_4779_inner <- mkFlatten(0);
    Operation_IFC mod_4779 <- mkDebugOperation(mod_4779_inner, "mod_4779");
    Operation_IFC mod_4780_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4780 <- mkDebugOperation(mod_4780_inner, "mod_4780");
    Operation_IFC mod_4781_inner <- mkUnaryMap(1680, silu_tile);
    Operation_IFC mod_4781 <- mkDebugOperation(mod_4781_inner, "mod_4781");
    Operation_IFC mod_4782_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4782 <- mkDebugOperation(mod_4782_inner, "mod_4782");
    Operation_IFC mod_4783_inner <- mkBinaryMap(1552, matmul_t_tile);
    Operation_IFC mod_4783 <- mkDebugOperation(mod_4783_inner, "mod_4783");
    PMU_IFC mod_4784_bufferize <- mkPMU(2);
    Operation_IFC mod_4784_inner = mod_4784_bufferize.operation;
    Operation_IFC mod_4784 <- mkDebugOperation(mod_4784_inner, "mod_4784");
    Operation_IFC mod_4785_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4785 <- mkDebugOperation(mod_4785_inner, "mod_4785");
    Operation_IFC mod_4786_inner <- mkFlatten(1);
    Operation_IFC mod_4786 <- mkDebugOperation(mod_4786_inner, "mod_4786");
    Operation_IFC mod_4787_inner <- mkFlatten(0);
    Operation_IFC mod_4787 <- mkDebugOperation(mod_4787_inner, "mod_4787");
    PMU_IFC mod_4788_bufferize <- mkPMU(1);
    Operation_IFC mod_4788_inner = mod_4788_bufferize.operation;
    Operation_IFC mod_4788 <- mkDebugOperation(mod_4788_inner, "mod_4788");
    Operation_IFC mod_4789_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4789 <- mkDebugOperation(mod_4789_inner, "mod_4789");
    PMU_IFC mod_4790_bufferize <- mkPMU(2);
    Operation_IFC mod_4790_inner = mod_4790_bufferize.operation;
    Operation_IFC mod_4790 <- mkDebugOperation(mod_4790_inner, "mod_4790");
    Operation_IFC mod_4791_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4791 <- mkDebugOperation(mod_4791_inner, "mod_4791");
    Operation_IFC mod_4792_inner <- mkFlatten(1);
    Operation_IFC mod_4792 <- mkDebugOperation(mod_4792_inner, "mod_4792");
    Operation_IFC mod_4793_inner <- mkFlatten(0);
    Operation_IFC mod_4793 <- mkDebugOperation(mod_4793_inner, "mod_4793");
    Operation_IFC mod_4794_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4794 <- mkDebugOperation(mod_4794_inner, "mod_4794");
    Operation_IFC mod_4795_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4795 <- mkDebugOperation(mod_4795_inner, "mod_4795");
    PMU_IFC mod_4796_bufferize <- mkPMU(2);
    Operation_IFC mod_4796_inner = mod_4796_bufferize.operation;
    Operation_IFC mod_4796 <- mkDebugOperation(mod_4796_inner, "mod_4796");
    rule rule_6149;
        ChannelMessage t;
        t <- mod_4771.get(1);
        mod_4772.put(0, t);
    endrule
    rule rule_6150;
        ChannelMessage t;
        t <- mod_4791.get(0);
        mod_4790.put(1, t);
    endrule
    rule rule_6151;
        ChannelMessage t;
        t <- mod_4775.get(1);
        mod_4771.put(1, t);
    endrule
    rule rule_6152;
        ChannelMessage t;
        t <- mod_4762.get(0);
        mod_4795.put(0, t);
    endrule
    rule rule_6153;
        ChannelMessage t;
        t <- mod_4762.get(1);
        mod_4763.put(0, t);
    endrule
    rule rule_6154;
        ChannelMessage t;
        t <- mod_4767.get(0);
        mod_4768.put(0, t);
    endrule
    rule rule_6155;
        ChannelMessage t;
        t <- mod_4795.get(0);
        mod_4762.put(1, t);
    endrule
    rule rule_6156;
        ChannelMessage t;
        t <- mod_4785.get(0);
        mod_4784.put(1, t);
    endrule
    rule rule_6157;
        ChannelMessage t;
        t <- mod_4768.get(0);
        mod_4780.put(0, t);
    endrule
    rule rule_6158;
        ChannelMessage t;
        t <- mod_4758.get(0);
        mod_4759.put(0, t);
    endrule
    rule rule_6159;
        ChannelMessage t;
        t <- mod_4775.get(0);
        mod_4775.put(1, t);
    endrule
    rule rule_6160;
        ChannelMessage t;
        t <- mod_4763.get(0);
        mod_4788.put(0, t);
    endrule
    rule rule_6161;
        ChannelMessage t;
        t <- mod_4796.get(1);
        mod_4760.put(1, t);
    endrule
    rule rule_6162;
        ChannelMessage t;
        t <- mod_4776.get(0);
        mod_4777.put(0, t);
    endrule
    rule rule_6163;
        ChannelMessage t;
        t <- mod_4786.get(0);
        mod_4784.put(0, t);
    endrule
    rule rule_6164;
        ChannelMessage t;
        t <- mod_4792.get(0);
        mod_4790.put(0, t);
    endrule
    rule rule_6165;
        ChannelMessage t;
        t <- mod_4794.get(0);
        mod_4764.put(1, t);
    endrule
    rule rule_6166;
        ChannelMessage t;
        t <- mod_4796.get(0);
        mod_4796.put(1, t);
    endrule
    rule rule_6167;
        ChannelMessage t;
        t <- mod_4787.get(0);
        mod_4786.put(0, t);
    endrule
    rule rule_6168;
        ChannelMessage t;
        t <- mod_4784.get(1);
        mod_4783.put(1, t);
    endrule
    rule rule_6169;
        ChannelMessage t;
        t <- mod_4765.get(0);
        mod_4766.put(0, t);
    endrule
    rule rule_6170;
        ChannelMessage t;
        t <- mod_4793.get(0);
        mod_4792.put(0, t);
    endrule
    rule rule_6171;
        ChannelMessage t;
        t <- mod_4788.get(0);
        mod_4789.put(0, t);
    endrule
    rule rule_6172;
        ChannelMessage t;
        t <- mod_4766.get(0);
        mod_4767.put(0, t);
    endrule
    rule rule_6173;
        ChannelMessage t;
        t <- mod_4760.get(0);
        mod_4796.put(0, t);
    endrule
    rule rule_6174;
        ChannelMessage t;
        t <- mod_4761.get(3);
        mod_4762.put(0, t);
    endrule
    rule rule_6175;
        ChannelMessage t;
        t <- mod_4757.get(0);
        mod_4758.put(0, t);
    endrule
    rule rule_6176;
        ChannelMessage t;
        t <- mod_4764.get(1);
        mod_4765.put(0, t);
    endrule
    rule rule_6177;
        ChannelMessage t;
        t <- mod_4781.get(0);
        mod_4767.put(1, t);
    endrule
    rule rule_6178;
        ChannelMessage t;
        t <- mod_4779.get(0);
        mod_4778.put(0, t);
    endrule
    rule rule_6179;
        ChannelMessage t;
        t <- mod_4768.get(1);
        mod_4769.put(0, t);
    endrule
    rule rule_6180;
        ChannelMessage t;
        t <- mod_4772.get(1);
        mod_4773.put(1, t);
    endrule
    rule rule_6181;
        ChannelMessage t;
        t <- mod_4774.get(0);
        mod_4774.put(1, t);
    endrule
    rule rule_6182;
        ChannelMessage t;
        t <- mod_4789.get(0);
        mod_4788.put(1, t);
    endrule
    rule rule_6183;
        ChannelMessage t;
        t <- mod_4778.get(0);
        mod_4776.put(0, t);
    endrule
    rule rule_6184;
        ChannelMessage t;
        t <- mod_4788.get(1);
        mod_4783.put(0, t);
    endrule
    rule rule_6185;
        ChannelMessage t;
        t <- mod_4760.get(1);
        mod_4761.put(0, t);
    endrule
    rule rule_6186;
        ChannelMessage t;
        t <- mod_4759.get(0);
        mod_4760.put(0, t);
    endrule
    rule rule_6187;
        ChannelMessage t;
        t <- mod_4774.get(1);
        mod_4772.put(1, t);
    endrule
    rule rule_6188;
        ChannelMessage t;
        t <- mod_4777.get(0);
        mod_4776.put(1, t);
    endrule
    rule rule_6189;
        ChannelMessage t;
        t <- mod_4770.get(0);
        mod_4771.put(0, t);
    endrule
    rule rule_6190;
        ChannelMessage t;
        t <- mod_4790.get(0);
        mod_4791.put(0, t);
    endrule
    rule rule_6191;
        ChannelMessage t;
        t <- mod_4769.get(0);
        mod_4770.put(0, t);
    endrule
    rule rule_6192;
        ChannelMessage t;
        t <- mod_4780.get(0);
        mod_4768.put(1, t);
    endrule
    rule rule_6193;
        ChannelMessage t;
        t <- mod_4771.get(0);
        mod_4775.put(0, t);
    endrule
    rule rule_6194;
        ChannelMessage t;
        t <- mod_4783.get(0);
        mod_4782.put(0, t);
    endrule
    rule rule_6195;
        ChannelMessage t;
        t <- mod_4790.get(1);
        mod_4765.put(1, t);
    endrule
    rule rule_6196;
        ChannelMessage t;
        t <- mod_4764.get(0);
        mod_4794.put(0, t);
    endrule
    rule rule_6197;
        ChannelMessage t;
        t <- mod_4784.get(0);
        mod_4785.put(0, t);
    endrule
    rule rule_6198;
        ChannelMessage t;
        t <- mod_4772.get(0);
        mod_4774.put(0, t);
    endrule
    rule rule_6199;
        ChannelMessage t;
        t <- mod_4763.get(1);
        mod_4764.put(0, t);
    endrule
    rule rule_6200;
        ChannelMessage t;
        t <- mod_4776.get(1);
        mod_4769.put(1, t);
    endrule
    rule rule_6201;
        ChannelMessage t;
        t <- mod_4782.get(0);
        mod_4781.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4757.put(0, t);
        end
        if (i == 1) begin
            mod_4773.put(0, t);
        end
        if (i == 2) begin
            mod_4779.put(0, t);
        end
        if (i == 3) begin
            mod_4787.put(0, t);
        end
        if (i == 4) begin
            mod_4793.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_4761.get(0);
        end
        if (i == 0) begin
            t <- mod_4761.get(1);
        end
        if (i == 2) begin
            t <- mod_4761.get(2);
        end
        if (i == 1) begin
            t <- mod_4773.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6151 (Operation_IFC);
    Operation_IFC mod_4798_inner <- mkReshape(2, 64);
    Operation_IFC mod_4798 <- mkDebugOperation(mod_4798_inner, "mod_4798");
    Operation_IFC mod_4799_inner <- mkFlatten(1);
    Operation_IFC mod_4799 <- mkDebugOperation(mod_4799_inner, "mod_4799");
    Operation_IFC mod_4800_inner <- mkFlatten(2);
    Operation_IFC mod_4800 <- mkDebugOperation(mod_4800_inner, "mod_4800");
    Operation_IFC mod_4801_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4801 <- mkDebugOperation(mod_4801_inner, "mod_4801");
    Broadcast_IFC#(4) mod_4802_inner <- mkBroadcast(4);
    Operation_IFC mod_4802 <- mkDebugOperation(mod_4802_inner.op, "mod_4802");
    PMU_IFC mod_4803_bufferize <- mkPMU(2);
    Operation_IFC mod_4803_inner = mod_4803_bufferize.operation;
    Operation_IFC mod_4803 <- mkDebugOperation(mod_4803_inner, "mod_4803");
    Broadcast_IFC#(2) mod_4804_inner <- mkBroadcast(2);
    Operation_IFC mod_4804 <- mkDebugOperation(mod_4804_inner.op, "mod_4804");
    PMU_IFC mod_4805_bufferize <- mkPMU(1);
    Operation_IFC mod_4805_inner = mod_4805_bufferize.operation;
    Operation_IFC mod_4805 <- mkDebugOperation(mod_4805_inner, "mod_4805");
    Operation_IFC mod_4806_inner <- mkBinaryMap(1039, matmul_t_tile);
    Operation_IFC mod_4806 <- mkDebugOperation(mod_4806_inner, "mod_4806");
    Operation_IFC mod_4807_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4807 <- mkDebugOperation(mod_4807_inner, "mod_4807");
    Operation_IFC mod_4808_inner <- mkBinaryMap(1807, mul_tile);
    Operation_IFC mod_4808 <- mkDebugOperation(mod_4808_inner, "mod_4808");
    PMU_IFC mod_4809_bufferize <- mkPMU(1);
    Operation_IFC mod_4809_inner = mod_4809_bufferize.operation;
    Operation_IFC mod_4809 <- mkDebugOperation(mod_4809_inner, "mod_4809");
    Operation_IFC mod_4810_inner <- mkBinaryMap(2329, matmul_t_tile);
    Operation_IFC mod_4810 <- mkDebugOperation(mod_4810_inner, "mod_4810");
    Operation_IFC mod_4811_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4811 <- mkDebugOperation(mod_4811_inner, "mod_4811");
    Operation_IFC mod_4812_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4812 <- mkDebugOperation(mod_4812_inner, "mod_4812");
    Operation_IFC mod_4813_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4813 <- mkDebugOperation(mod_4813_inner, "mod_4813");
    Operation_IFC mod_4814_inner <- mkBinaryMap(2706, mul_tile);
    Operation_IFC mod_4814 <- mkDebugOperation(mod_4814_inner, "mod_4814");
    PMU_IFC mod_4815_bufferize <- mkPMU(1);
    Operation_IFC mod_4815_inner = mod_4815_bufferize.operation;
    Operation_IFC mod_4815 <- mkDebugOperation(mod_4815_inner, "mod_4815");
    PMU_IFC mod_4816_bufferize <- mkPMU(2);
    Operation_IFC mod_4816_inner = mod_4816_bufferize.operation;
    Operation_IFC mod_4816 <- mkDebugOperation(mod_4816_inner, "mod_4816");
    PMU_IFC mod_4817_bufferize <- mkPMU(2);
    Operation_IFC mod_4817_inner = mod_4817_bufferize.operation;
    Operation_IFC mod_4817 <- mkDebugOperation(mod_4817_inner, "mod_4817");
    Operation_IFC mod_4818_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4818 <- mkDebugOperation(mod_4818_inner, "mod_4818");
    Operation_IFC mod_4819_inner <- mkFlatten(1);
    Operation_IFC mod_4819 <- mkDebugOperation(mod_4819_inner, "mod_4819");
    Operation_IFC mod_4820_inner <- mkFlatten(0);
    Operation_IFC mod_4820 <- mkDebugOperation(mod_4820_inner, "mod_4820");
    Operation_IFC mod_4821_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4821 <- mkDebugOperation(mod_4821_inner, "mod_4821");
    Operation_IFC mod_4822_inner <- mkUnaryMap(1679, silu_tile);
    Operation_IFC mod_4822 <- mkDebugOperation(mod_4822_inner, "mod_4822");
    Operation_IFC mod_4823_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4823 <- mkDebugOperation(mod_4823_inner, "mod_4823");
    Operation_IFC mod_4824_inner <- mkBinaryMap(1551, matmul_t_tile);
    Operation_IFC mod_4824 <- mkDebugOperation(mod_4824_inner, "mod_4824");
    PMU_IFC mod_4825_bufferize <- mkPMU(2);
    Operation_IFC mod_4825_inner = mod_4825_bufferize.operation;
    Operation_IFC mod_4825 <- mkDebugOperation(mod_4825_inner, "mod_4825");
    Operation_IFC mod_4826_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4826 <- mkDebugOperation(mod_4826_inner, "mod_4826");
    Operation_IFC mod_4827_inner <- mkFlatten(1);
    Operation_IFC mod_4827 <- mkDebugOperation(mod_4827_inner, "mod_4827");
    Operation_IFC mod_4828_inner <- mkFlatten(0);
    Operation_IFC mod_4828 <- mkDebugOperation(mod_4828_inner, "mod_4828");
    PMU_IFC mod_4829_bufferize <- mkPMU(1);
    Operation_IFC mod_4829_inner = mod_4829_bufferize.operation;
    Operation_IFC mod_4829 <- mkDebugOperation(mod_4829_inner, "mod_4829");
    Operation_IFC mod_4830_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4830 <- mkDebugOperation(mod_4830_inner, "mod_4830");
    PMU_IFC mod_4831_bufferize <- mkPMU(2);
    Operation_IFC mod_4831_inner = mod_4831_bufferize.operation;
    Operation_IFC mod_4831 <- mkDebugOperation(mod_4831_inner, "mod_4831");
    Operation_IFC mod_4832_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4832 <- mkDebugOperation(mod_4832_inner, "mod_4832");
    Operation_IFC mod_4833_inner <- mkFlatten(1);
    Operation_IFC mod_4833 <- mkDebugOperation(mod_4833_inner, "mod_4833");
    Operation_IFC mod_4834_inner <- mkFlatten(0);
    Operation_IFC mod_4834 <- mkDebugOperation(mod_4834_inner, "mod_4834");
    Operation_IFC mod_4835_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4835 <- mkDebugOperation(mod_4835_inner, "mod_4835");
    Operation_IFC mod_4836_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4836 <- mkDebugOperation(mod_4836_inner, "mod_4836");
    PMU_IFC mod_4837_bufferize <- mkPMU(2);
    Operation_IFC mod_4837_inner = mod_4837_bufferize.operation;
    Operation_IFC mod_4837 <- mkDebugOperation(mod_4837_inner, "mod_4837");
    rule rule_6202;
        ChannelMessage t;
        t <- mod_4835.get(0);
        mod_4805.put(1, t);
    endrule
    rule rule_6203;
        ChannelMessage t;
        t <- mod_4815.get(1);
        mod_4813.put(1, t);
    endrule
    rule rule_6204;
        ChannelMessage t;
        t <- mod_4818.get(0);
        mod_4817.put(1, t);
    endrule
    rule rule_6205;
        ChannelMessage t;
        t <- mod_4815.get(0);
        mod_4815.put(1, t);
    endrule
    rule rule_6206;
        ChannelMessage t;
        t <- mod_4831.get(0);
        mod_4832.put(0, t);
    endrule
    rule rule_6207;
        ChannelMessage t;
        t <- mod_4810.get(0);
        mod_4811.put(0, t);
    endrule
    rule rule_6208;
        ChannelMessage t;
        t <- mod_4813.get(0);
        mod_4815.put(0, t);
    endrule
    rule rule_6209;
        ChannelMessage t;
        t <- mod_4819.get(0);
        mod_4817.put(0, t);
    endrule
    rule rule_6210;
        ChannelMessage t;
        t <- mod_4816.get(0);
        mod_4816.put(1, t);
    endrule
    rule rule_6211;
        ChannelMessage t;
        t <- mod_4832.get(0);
        mod_4831.put(1, t);
    endrule
    rule rule_6212;
        ChannelMessage t;
        t <- mod_4817.get(0);
        mod_4818.put(0, t);
    endrule
    rule rule_6213;
        ChannelMessage t;
        t <- mod_4834.get(0);
        mod_4833.put(0, t);
    endrule
    rule rule_6214;
        ChannelMessage t;
        t <- mod_4812.get(1);
        mod_4813.put(0, t);
    endrule
    rule rule_6215;
        ChannelMessage t;
        t <- mod_4820.get(0);
        mod_4819.put(0, t);
    endrule
    rule rule_6216;
        ChannelMessage t;
        t <- mod_4821.get(0);
        mod_4809.put(1, t);
    endrule
    rule rule_6217;
        ChannelMessage t;
        t <- mod_4802.get(3);
        mod_4803.put(0, t);
    endrule
    rule rule_6218;
        ChannelMessage t;
        t <- mod_4837.get(1);
        mod_4801.put(1, t);
    endrule
    rule rule_6219;
        ChannelMessage t;
        t <- mod_4813.get(1);
        mod_4814.put(1, t);
    endrule
    rule rule_6220;
        ChannelMessage t;
        t <- mod_4807.get(0);
        mod_4808.put(0, t);
    endrule
    rule rule_6221;
        ChannelMessage t;
        t <- mod_4817.get(1);
        mod_4810.put(1, t);
    endrule
    rule rule_6222;
        ChannelMessage t;
        t <- mod_4803.get(0);
        mod_4836.put(0, t);
    endrule
    rule rule_6223;
        ChannelMessage t;
        t <- mod_4809.get(0);
        mod_4821.put(0, t);
    endrule
    rule rule_6224;
        ChannelMessage t;
        t <- mod_4808.get(0);
        mod_4809.put(0, t);
    endrule
    rule rule_6225;
        ChannelMessage t;
        t <- mod_4831.get(1);
        mod_4806.put(1, t);
    endrule
    rule rule_6226;
        ChannelMessage t;
        t <- mod_4798.get(0);
        mod_4799.put(0, t);
    endrule
    rule rule_6227;
        ChannelMessage t;
        t <- mod_4804.get(1);
        mod_4805.put(0, t);
    endrule
    rule rule_6228;
        ChannelMessage t;
        t <- mod_4806.get(0);
        mod_4807.put(0, t);
    endrule
    rule rule_6229;
        ChannelMessage t;
        t <- mod_4837.get(0);
        mod_4837.put(1, t);
    endrule
    rule rule_6230;
        ChannelMessage t;
        t <- mod_4824.get(0);
        mod_4823.put(0, t);
    endrule
    rule rule_6231;
        ChannelMessage t;
        t <- mod_4799.get(0);
        mod_4800.put(0, t);
    endrule
    rule rule_6232;
        ChannelMessage t;
        t <- mod_4830.get(0);
        mod_4829.put(1, t);
    endrule
    rule rule_6233;
        ChannelMessage t;
        t <- mod_4816.get(1);
        mod_4812.put(1, t);
    endrule
    rule rule_6234;
        ChannelMessage t;
        t <- mod_4803.get(1);
        mod_4804.put(0, t);
    endrule
    rule rule_6235;
        ChannelMessage t;
        t <- mod_4801.get(0);
        mod_4837.put(0, t);
    endrule
    rule rule_6236;
        ChannelMessage t;
        t <- mod_4836.get(0);
        mod_4803.put(1, t);
    endrule
    rule rule_6237;
        ChannelMessage t;
        t <- mod_4825.get(0);
        mod_4826.put(0, t);
    endrule
    rule rule_6238;
        ChannelMessage t;
        t <- mod_4826.get(0);
        mod_4825.put(1, t);
    endrule
    rule rule_6239;
        ChannelMessage t;
        t <- mod_4822.get(0);
        mod_4808.put(1, t);
    endrule
    rule rule_6240;
        ChannelMessage t;
        t <- mod_4829.get(0);
        mod_4830.put(0, t);
    endrule
    rule rule_6241;
        ChannelMessage t;
        t <- mod_4800.get(0);
        mod_4801.put(0, t);
    endrule
    rule rule_6242;
        ChannelMessage t;
        t <- mod_4829.get(1);
        mod_4824.put(0, t);
    endrule
    rule rule_6243;
        ChannelMessage t;
        t <- mod_4801.get(1);
        mod_4802.put(0, t);
    endrule
    rule rule_6244;
        ChannelMessage t;
        t <- mod_4833.get(0);
        mod_4831.put(0, t);
    endrule
    rule rule_6245;
        ChannelMessage t;
        t <- mod_4827.get(0);
        mod_4825.put(0, t);
    endrule
    rule rule_6246;
        ChannelMessage t;
        t <- mod_4811.get(0);
        mod_4812.put(0, t);
    endrule
    rule rule_6247;
        ChannelMessage t;
        t <- mod_4825.get(1);
        mod_4824.put(1, t);
    endrule
    rule rule_6248;
        ChannelMessage t;
        t <- mod_4805.get(1);
        mod_4806.put(0, t);
    endrule
    rule rule_6249;
        ChannelMessage t;
        t <- mod_4804.get(0);
        mod_4829.put(0, t);
    endrule
    rule rule_6250;
        ChannelMessage t;
        t <- mod_4809.get(1);
        mod_4810.put(0, t);
    endrule
    rule rule_6251;
        ChannelMessage t;
        t <- mod_4812.get(0);
        mod_4816.put(0, t);
    endrule
    rule rule_6252;
        ChannelMessage t;
        t <- mod_4805.get(0);
        mod_4835.put(0, t);
    endrule
    rule rule_6253;
        ChannelMessage t;
        t <- mod_4823.get(0);
        mod_4822.put(0, t);
    endrule
    rule rule_6254;
        ChannelMessage t;
        t <- mod_4828.get(0);
        mod_4827.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4798.put(0, t);
        end
        if (i == 1) begin
            mod_4814.put(0, t);
        end
        if (i == 2) begin
            mod_4820.put(0, t);
        end
        if (i == 3) begin
            mod_4828.put(0, t);
        end
        if (i == 4) begin
            mod_4834.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 2) begin
            t <- mod_4802.get(0);
        end
        if (i == 0) begin
            t <- mod_4802.get(1);
        end
        if (i == 1) begin
            t <- mod_4802.get(2);
        end
        if (i == 3) begin
            t <- mod_4814.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6152 (Operation_IFC);
    Operation_IFC mod_4839_inner <- mkReshape(2, 64);
    Operation_IFC mod_4839 <- mkDebugOperation(mod_4839_inner, "mod_4839");
    Operation_IFC mod_4840_inner <- mkFlatten(1);
    Operation_IFC mod_4840 <- mkDebugOperation(mod_4840_inner, "mod_4840");
    Operation_IFC mod_4841_inner <- mkFlatten(2);
    Operation_IFC mod_4841 <- mkDebugOperation(mod_4841_inner, "mod_4841");
    Operation_IFC mod_4842_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4842 <- mkDebugOperation(mod_4842_inner, "mod_4842");
    Broadcast_IFC#(4) mod_4843_inner <- mkBroadcast(4);
    Operation_IFC mod_4843 <- mkDebugOperation(mod_4843_inner.op, "mod_4843");
    PMU_IFC mod_4844_bufferize <- mkPMU(2);
    Operation_IFC mod_4844_inner = mod_4844_bufferize.operation;
    Operation_IFC mod_4844 <- mkDebugOperation(mod_4844_inner, "mod_4844");
    Broadcast_IFC#(2) mod_4845_inner <- mkBroadcast(2);
    Operation_IFC mod_4845 <- mkDebugOperation(mod_4845_inner.op, "mod_4845");
    PMU_IFC mod_4846_bufferize <- mkPMU(1);
    Operation_IFC mod_4846_inner = mod_4846_bufferize.operation;
    Operation_IFC mod_4846 <- mkDebugOperation(mod_4846_inner, "mod_4846");
    Operation_IFC mod_4847_inner <- mkBinaryMap(1038, matmul_t_tile);
    Operation_IFC mod_4847 <- mkDebugOperation(mod_4847_inner, "mod_4847");
    Operation_IFC mod_4848_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4848 <- mkDebugOperation(mod_4848_inner, "mod_4848");
    Operation_IFC mod_4849_inner <- mkBinaryMap(1806, mul_tile);
    Operation_IFC mod_4849 <- mkDebugOperation(mod_4849_inner, "mod_4849");
    PMU_IFC mod_4850_bufferize <- mkPMU(1);
    Operation_IFC mod_4850_inner = mod_4850_bufferize.operation;
    Operation_IFC mod_4850 <- mkDebugOperation(mod_4850_inner, "mod_4850");
    Operation_IFC mod_4851_inner <- mkBinaryMap(2327, matmul_t_tile);
    Operation_IFC mod_4851 <- mkDebugOperation(mod_4851_inner, "mod_4851");
    Operation_IFC mod_4852_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4852 <- mkDebugOperation(mod_4852_inner, "mod_4852");
    Operation_IFC mod_4853_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4853 <- mkDebugOperation(mod_4853_inner, "mod_4853");
    Operation_IFC mod_4854_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4854 <- mkDebugOperation(mod_4854_inner, "mod_4854");
    Operation_IFC mod_4855_inner <- mkBinaryMap(2705, mul_tile);
    Operation_IFC mod_4855 <- mkDebugOperation(mod_4855_inner, "mod_4855");
    PMU_IFC mod_4856_bufferize <- mkPMU(1);
    Operation_IFC mod_4856_inner = mod_4856_bufferize.operation;
    Operation_IFC mod_4856 <- mkDebugOperation(mod_4856_inner, "mod_4856");
    PMU_IFC mod_4857_bufferize <- mkPMU(2);
    Operation_IFC mod_4857_inner = mod_4857_bufferize.operation;
    Operation_IFC mod_4857 <- mkDebugOperation(mod_4857_inner, "mod_4857");
    PMU_IFC mod_4858_bufferize <- mkPMU(2);
    Operation_IFC mod_4858_inner = mod_4858_bufferize.operation;
    Operation_IFC mod_4858 <- mkDebugOperation(mod_4858_inner, "mod_4858");
    Operation_IFC mod_4859_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4859 <- mkDebugOperation(mod_4859_inner, "mod_4859");
    Operation_IFC mod_4860_inner <- mkFlatten(1);
    Operation_IFC mod_4860 <- mkDebugOperation(mod_4860_inner, "mod_4860");
    Operation_IFC mod_4861_inner <- mkFlatten(0);
    Operation_IFC mod_4861 <- mkDebugOperation(mod_4861_inner, "mod_4861");
    Operation_IFC mod_4862_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4862 <- mkDebugOperation(mod_4862_inner, "mod_4862");
    Operation_IFC mod_4863_inner <- mkUnaryMap(1678, silu_tile);
    Operation_IFC mod_4863 <- mkDebugOperation(mod_4863_inner, "mod_4863");
    Operation_IFC mod_4864_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4864 <- mkDebugOperation(mod_4864_inner, "mod_4864");
    Operation_IFC mod_4865_inner <- mkBinaryMap(1550, matmul_t_tile);
    Operation_IFC mod_4865 <- mkDebugOperation(mod_4865_inner, "mod_4865");
    PMU_IFC mod_4866_bufferize <- mkPMU(2);
    Operation_IFC mod_4866_inner = mod_4866_bufferize.operation;
    Operation_IFC mod_4866 <- mkDebugOperation(mod_4866_inner, "mod_4866");
    Operation_IFC mod_4867_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4867 <- mkDebugOperation(mod_4867_inner, "mod_4867");
    Operation_IFC mod_4868_inner <- mkFlatten(1);
    Operation_IFC mod_4868 <- mkDebugOperation(mod_4868_inner, "mod_4868");
    Operation_IFC mod_4869_inner <- mkFlatten(0);
    Operation_IFC mod_4869 <- mkDebugOperation(mod_4869_inner, "mod_4869");
    PMU_IFC mod_4870_bufferize <- mkPMU(1);
    Operation_IFC mod_4870_inner = mod_4870_bufferize.operation;
    Operation_IFC mod_4870 <- mkDebugOperation(mod_4870_inner, "mod_4870");
    Operation_IFC mod_4871_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4871 <- mkDebugOperation(mod_4871_inner, "mod_4871");
    PMU_IFC mod_4872_bufferize <- mkPMU(2);
    Operation_IFC mod_4872_inner = mod_4872_bufferize.operation;
    Operation_IFC mod_4872 <- mkDebugOperation(mod_4872_inner, "mod_4872");
    Operation_IFC mod_4873_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4873 <- mkDebugOperation(mod_4873_inner, "mod_4873");
    Operation_IFC mod_4874_inner <- mkFlatten(1);
    Operation_IFC mod_4874 <- mkDebugOperation(mod_4874_inner, "mod_4874");
    Operation_IFC mod_4875_inner <- mkFlatten(0);
    Operation_IFC mod_4875 <- mkDebugOperation(mod_4875_inner, "mod_4875");
    Operation_IFC mod_4876_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4876 <- mkDebugOperation(mod_4876_inner, "mod_4876");
    Operation_IFC mod_4877_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4877 <- mkDebugOperation(mod_4877_inner, "mod_4877");
    PMU_IFC mod_4878_bufferize <- mkPMU(2);
    Operation_IFC mod_4878_inner = mod_4878_bufferize.operation;
    Operation_IFC mod_4878 <- mkDebugOperation(mod_4878_inner, "mod_4878");
    rule rule_6255;
        ChannelMessage t;
        t <- mod_4861.get(0);
        mod_4860.put(0, t);
    endrule
    rule rule_6256;
        ChannelMessage t;
        t <- mod_4856.get(1);
        mod_4854.put(1, t);
    endrule
    rule rule_6257;
        ChannelMessage t;
        t <- mod_4849.get(0);
        mod_4850.put(0, t);
    endrule
    rule rule_6258;
        ChannelMessage t;
        t <- mod_4843.get(3);
        mod_4844.put(0, t);
    endrule
    rule rule_6259;
        ChannelMessage t;
        t <- mod_4844.get(1);
        mod_4845.put(0, t);
    endrule
    rule rule_6260;
        ChannelMessage t;
        t <- mod_4859.get(0);
        mod_4858.put(1, t);
    endrule
    rule rule_6261;
        ChannelMessage t;
        t <- mod_4840.get(0);
        mod_4841.put(0, t);
    endrule
    rule rule_6262;
        ChannelMessage t;
        t <- mod_4870.get(0);
        mod_4871.put(0, t);
    endrule
    rule rule_6263;
        ChannelMessage t;
        t <- mod_4873.get(0);
        mod_4872.put(1, t);
    endrule
    rule rule_6264;
        ChannelMessage t;
        t <- mod_4853.get(1);
        mod_4854.put(0, t);
    endrule
    rule rule_6265;
        ChannelMessage t;
        t <- mod_4864.get(0);
        mod_4863.put(0, t);
    endrule
    rule rule_6266;
        ChannelMessage t;
        t <- mod_4853.get(0);
        mod_4857.put(0, t);
    endrule
    rule rule_6267;
        ChannelMessage t;
        t <- mod_4857.get(0);
        mod_4857.put(1, t);
    endrule
    rule rule_6268;
        ChannelMessage t;
        t <- mod_4870.get(1);
        mod_4865.put(0, t);
    endrule
    rule rule_6269;
        ChannelMessage t;
        t <- mod_4871.get(0);
        mod_4870.put(1, t);
    endrule
    rule rule_6270;
        ChannelMessage t;
        t <- mod_4866.get(0);
        mod_4867.put(0, t);
    endrule
    rule rule_6271;
        ChannelMessage t;
        t <- mod_4872.get(0);
        mod_4873.put(0, t);
    endrule
    rule rule_6272;
        ChannelMessage t;
        t <- mod_4850.get(0);
        mod_4862.put(0, t);
    endrule
    rule rule_6273;
        ChannelMessage t;
        t <- mod_4878.get(1);
        mod_4842.put(1, t);
    endrule
    rule rule_6274;
        ChannelMessage t;
        t <- mod_4872.get(1);
        mod_4847.put(1, t);
    endrule
    rule rule_6275;
        ChannelMessage t;
        t <- mod_4875.get(0);
        mod_4874.put(0, t);
    endrule
    rule rule_6276;
        ChannelMessage t;
        t <- mod_4842.get(1);
        mod_4843.put(0, t);
    endrule
    rule rule_6277;
        ChannelMessage t;
        t <- mod_4867.get(0);
        mod_4866.put(1, t);
    endrule
    rule rule_6278;
        ChannelMessage t;
        t <- mod_4878.get(0);
        mod_4878.put(1, t);
    endrule
    rule rule_6279;
        ChannelMessage t;
        t <- mod_4851.get(0);
        mod_4852.put(0, t);
    endrule
    rule rule_6280;
        ChannelMessage t;
        t <- mod_4848.get(0);
        mod_4849.put(0, t);
    endrule
    rule rule_6281;
        ChannelMessage t;
        t <- mod_4850.get(1);
        mod_4851.put(0, t);
    endrule
    rule rule_6282;
        ChannelMessage t;
        t <- mod_4857.get(1);
        mod_4853.put(1, t);
    endrule
    rule rule_6283;
        ChannelMessage t;
        t <- mod_4852.get(0);
        mod_4853.put(0, t);
    endrule
    rule rule_6284;
        ChannelMessage t;
        t <- mod_4842.get(0);
        mod_4878.put(0, t);
    endrule
    rule rule_6285;
        ChannelMessage t;
        t <- mod_4854.get(0);
        mod_4856.put(0, t);
    endrule
    rule rule_6286;
        ChannelMessage t;
        t <- mod_4858.get(1);
        mod_4851.put(1, t);
    endrule
    rule rule_6287;
        ChannelMessage t;
        t <- mod_4868.get(0);
        mod_4866.put(0, t);
    endrule
    rule rule_6288;
        ChannelMessage t;
        t <- mod_4863.get(0);
        mod_4849.put(1, t);
    endrule
    rule rule_6289;
        ChannelMessage t;
        t <- mod_4869.get(0);
        mod_4868.put(0, t);
    endrule
    rule rule_6290;
        ChannelMessage t;
        t <- mod_4839.get(0);
        mod_4840.put(0, t);
    endrule
    rule rule_6291;
        ChannelMessage t;
        t <- mod_4876.get(0);
        mod_4846.put(1, t);
    endrule
    rule rule_6292;
        ChannelMessage t;
        t <- mod_4854.get(1);
        mod_4855.put(1, t);
    endrule
    rule rule_6293;
        ChannelMessage t;
        t <- mod_4874.get(0);
        mod_4872.put(0, t);
    endrule
    rule rule_6294;
        ChannelMessage t;
        t <- mod_4846.get(1);
        mod_4847.put(0, t);
    endrule
    rule rule_6295;
        ChannelMessage t;
        t <- mod_4847.get(0);
        mod_4848.put(0, t);
    endrule
    rule rule_6296;
        ChannelMessage t;
        t <- mod_4860.get(0);
        mod_4858.put(0, t);
    endrule
    rule rule_6297;
        ChannelMessage t;
        t <- mod_4865.get(0);
        mod_4864.put(0, t);
    endrule
    rule rule_6298;
        ChannelMessage t;
        t <- mod_4846.get(0);
        mod_4876.put(0, t);
    endrule
    rule rule_6299;
        ChannelMessage t;
        t <- mod_4844.get(0);
        mod_4877.put(0, t);
    endrule
    rule rule_6300;
        ChannelMessage t;
        t <- mod_4845.get(1);
        mod_4846.put(0, t);
    endrule
    rule rule_6301;
        ChannelMessage t;
        t <- mod_4845.get(0);
        mod_4870.put(0, t);
    endrule
    rule rule_6302;
        ChannelMessage t;
        t <- mod_4858.get(0);
        mod_4859.put(0, t);
    endrule
    rule rule_6303;
        ChannelMessage t;
        t <- mod_4877.get(0);
        mod_4844.put(1, t);
    endrule
    rule rule_6304;
        ChannelMessage t;
        t <- mod_4862.get(0);
        mod_4850.put(1, t);
    endrule
    rule rule_6305;
        ChannelMessage t;
        t <- mod_4856.get(0);
        mod_4856.put(1, t);
    endrule
    rule rule_6306;
        ChannelMessage t;
        t <- mod_4866.get(1);
        mod_4865.put(1, t);
    endrule
    rule rule_6307;
        ChannelMessage t;
        t <- mod_4841.get(0);
        mod_4842.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4839.put(0, t);
        end
        if (i == 1) begin
            mod_4855.put(0, t);
        end
        if (i == 2) begin
            mod_4861.put(0, t);
        end
        if (i == 3) begin
            mod_4869.put(0, t);
        end
        if (i == 4) begin
            mod_4875.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_4843.get(0);
        end
        if (i == 0) begin
            t <- mod_4843.get(1);
        end
        if (i == 3) begin
            t <- mod_4843.get(2);
        end
        if (i == 2) begin
            t <- mod_4855.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6153 (Operation_IFC);
    Operation_IFC mod_4880_inner <- mkReshape(2, 64);
    Operation_IFC mod_4880 <- mkDebugOperation(mod_4880_inner, "mod_4880");
    Operation_IFC mod_4881_inner <- mkFlatten(1);
    Operation_IFC mod_4881 <- mkDebugOperation(mod_4881_inner, "mod_4881");
    Operation_IFC mod_4882_inner <- mkFlatten(2);
    Operation_IFC mod_4882 <- mkDebugOperation(mod_4882_inner, "mod_4882");
    Operation_IFC mod_4883_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4883 <- mkDebugOperation(mod_4883_inner, "mod_4883");
    Broadcast_IFC#(4) mod_4884_inner <- mkBroadcast(4);
    Operation_IFC mod_4884 <- mkDebugOperation(mod_4884_inner.op, "mod_4884");
    PMU_IFC mod_4885_bufferize <- mkPMU(2);
    Operation_IFC mod_4885_inner = mod_4885_bufferize.operation;
    Operation_IFC mod_4885 <- mkDebugOperation(mod_4885_inner, "mod_4885");
    Broadcast_IFC#(2) mod_4886_inner <- mkBroadcast(2);
    Operation_IFC mod_4886 <- mkDebugOperation(mod_4886_inner.op, "mod_4886");
    PMU_IFC mod_4887_bufferize <- mkPMU(1);
    Operation_IFC mod_4887_inner = mod_4887_bufferize.operation;
    Operation_IFC mod_4887 <- mkDebugOperation(mod_4887_inner, "mod_4887");
    Operation_IFC mod_4888_inner <- mkBinaryMap(1037, matmul_t_tile);
    Operation_IFC mod_4888 <- mkDebugOperation(mod_4888_inner, "mod_4888");
    Operation_IFC mod_4889_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4889 <- mkDebugOperation(mod_4889_inner, "mod_4889");
    Operation_IFC mod_4890_inner <- mkBinaryMap(1805, mul_tile);
    Operation_IFC mod_4890 <- mkDebugOperation(mod_4890_inner, "mod_4890");
    PMU_IFC mod_4891_bufferize <- mkPMU(1);
    Operation_IFC mod_4891_inner = mod_4891_bufferize.operation;
    Operation_IFC mod_4891 <- mkDebugOperation(mod_4891_inner, "mod_4891");
    Operation_IFC mod_4892_inner <- mkBinaryMap(2325, matmul_t_tile);
    Operation_IFC mod_4892 <- mkDebugOperation(mod_4892_inner, "mod_4892");
    Operation_IFC mod_4893_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4893 <- mkDebugOperation(mod_4893_inner, "mod_4893");
    Operation_IFC mod_4894_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4894 <- mkDebugOperation(mod_4894_inner, "mod_4894");
    Operation_IFC mod_4895_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4895 <- mkDebugOperation(mod_4895_inner, "mod_4895");
    Operation_IFC mod_4896_inner <- mkBinaryMap(2704, mul_tile);
    Operation_IFC mod_4896 <- mkDebugOperation(mod_4896_inner, "mod_4896");
    PMU_IFC mod_4897_bufferize <- mkPMU(1);
    Operation_IFC mod_4897_inner = mod_4897_bufferize.operation;
    Operation_IFC mod_4897 <- mkDebugOperation(mod_4897_inner, "mod_4897");
    PMU_IFC mod_4898_bufferize <- mkPMU(2);
    Operation_IFC mod_4898_inner = mod_4898_bufferize.operation;
    Operation_IFC mod_4898 <- mkDebugOperation(mod_4898_inner, "mod_4898");
    PMU_IFC mod_4899_bufferize <- mkPMU(2);
    Operation_IFC mod_4899_inner = mod_4899_bufferize.operation;
    Operation_IFC mod_4899 <- mkDebugOperation(mod_4899_inner, "mod_4899");
    Operation_IFC mod_4900_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4900 <- mkDebugOperation(mod_4900_inner, "mod_4900");
    Operation_IFC mod_4901_inner <- mkFlatten(1);
    Operation_IFC mod_4901 <- mkDebugOperation(mod_4901_inner, "mod_4901");
    Operation_IFC mod_4902_inner <- mkFlatten(0);
    Operation_IFC mod_4902 <- mkDebugOperation(mod_4902_inner, "mod_4902");
    Operation_IFC mod_4903_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4903 <- mkDebugOperation(mod_4903_inner, "mod_4903");
    Operation_IFC mod_4904_inner <- mkUnaryMap(1677, silu_tile);
    Operation_IFC mod_4904 <- mkDebugOperation(mod_4904_inner, "mod_4904");
    Operation_IFC mod_4905_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4905 <- mkDebugOperation(mod_4905_inner, "mod_4905");
    Operation_IFC mod_4906_inner <- mkBinaryMap(1549, matmul_t_tile);
    Operation_IFC mod_4906 <- mkDebugOperation(mod_4906_inner, "mod_4906");
    PMU_IFC mod_4907_bufferize <- mkPMU(2);
    Operation_IFC mod_4907_inner = mod_4907_bufferize.operation;
    Operation_IFC mod_4907 <- mkDebugOperation(mod_4907_inner, "mod_4907");
    Operation_IFC mod_4908_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4908 <- mkDebugOperation(mod_4908_inner, "mod_4908");
    Operation_IFC mod_4909_inner <- mkFlatten(1);
    Operation_IFC mod_4909 <- mkDebugOperation(mod_4909_inner, "mod_4909");
    Operation_IFC mod_4910_inner <- mkFlatten(0);
    Operation_IFC mod_4910 <- mkDebugOperation(mod_4910_inner, "mod_4910");
    PMU_IFC mod_4911_bufferize <- mkPMU(1);
    Operation_IFC mod_4911_inner = mod_4911_bufferize.operation;
    Operation_IFC mod_4911 <- mkDebugOperation(mod_4911_inner, "mod_4911");
    Operation_IFC mod_4912_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4912 <- mkDebugOperation(mod_4912_inner, "mod_4912");
    PMU_IFC mod_4913_bufferize <- mkPMU(2);
    Operation_IFC mod_4913_inner = mod_4913_bufferize.operation;
    Operation_IFC mod_4913 <- mkDebugOperation(mod_4913_inner, "mod_4913");
    Operation_IFC mod_4914_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4914 <- mkDebugOperation(mod_4914_inner, "mod_4914");
    Operation_IFC mod_4915_inner <- mkFlatten(1);
    Operation_IFC mod_4915 <- mkDebugOperation(mod_4915_inner, "mod_4915");
    Operation_IFC mod_4916_inner <- mkFlatten(0);
    Operation_IFC mod_4916 <- mkDebugOperation(mod_4916_inner, "mod_4916");
    Operation_IFC mod_4917_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4917 <- mkDebugOperation(mod_4917_inner, "mod_4917");
    Operation_IFC mod_4918_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4918 <- mkDebugOperation(mod_4918_inner, "mod_4918");
    PMU_IFC mod_4919_bufferize <- mkPMU(2);
    Operation_IFC mod_4919_inner = mod_4919_bufferize.operation;
    Operation_IFC mod_4919 <- mkDebugOperation(mod_4919_inner, "mod_4919");
    rule rule_6308;
        ChannelMessage t;
        t <- mod_4891.get(0);
        mod_4903.put(0, t);
    endrule
    rule rule_6309;
        ChannelMessage t;
        t <- mod_4898.get(1);
        mod_4894.put(1, t);
    endrule
    rule rule_6310;
        ChannelMessage t;
        t <- mod_4895.get(1);
        mod_4896.put(1, t);
    endrule
    rule rule_6311;
        ChannelMessage t;
        t <- mod_4905.get(0);
        mod_4904.put(0, t);
    endrule
    rule rule_6312;
        ChannelMessage t;
        t <- mod_4903.get(0);
        mod_4891.put(1, t);
    endrule
    rule rule_6313;
        ChannelMessage t;
        t <- mod_4913.get(0);
        mod_4914.put(0, t);
    endrule
    rule rule_6314;
        ChannelMessage t;
        t <- mod_4917.get(0);
        mod_4887.put(1, t);
    endrule
    rule rule_6315;
        ChannelMessage t;
        t <- mod_4919.get(0);
        mod_4919.put(1, t);
    endrule
    rule rule_6316;
        ChannelMessage t;
        t <- mod_4880.get(0);
        mod_4881.put(0, t);
    endrule
    rule rule_6317;
        ChannelMessage t;
        t <- mod_4897.get(0);
        mod_4897.put(1, t);
    endrule
    rule rule_6318;
        ChannelMessage t;
        t <- mod_4916.get(0);
        mod_4915.put(0, t);
    endrule
    rule rule_6319;
        ChannelMessage t;
        t <- mod_4918.get(0);
        mod_4885.put(1, t);
    endrule
    rule rule_6320;
        ChannelMessage t;
        t <- mod_4894.get(1);
        mod_4895.put(0, t);
    endrule
    rule rule_6321;
        ChannelMessage t;
        t <- mod_4919.get(1);
        mod_4883.put(1, t);
    endrule
    rule rule_6322;
        ChannelMessage t;
        t <- mod_4885.get(1);
        mod_4886.put(0, t);
    endrule
    rule rule_6323;
        ChannelMessage t;
        t <- mod_4907.get(0);
        mod_4908.put(0, t);
    endrule
    rule rule_6324;
        ChannelMessage t;
        t <- mod_4886.get(1);
        mod_4887.put(0, t);
    endrule
    rule rule_6325;
        ChannelMessage t;
        t <- mod_4887.get(1);
        mod_4888.put(0, t);
    endrule
    rule rule_6326;
        ChannelMessage t;
        t <- mod_4901.get(0);
        mod_4899.put(0, t);
    endrule
    rule rule_6327;
        ChannelMessage t;
        t <- mod_4885.get(0);
        mod_4918.put(0, t);
    endrule
    rule rule_6328;
        ChannelMessage t;
        t <- mod_4894.get(0);
        mod_4898.put(0, t);
    endrule
    rule rule_6329;
        ChannelMessage t;
        t <- mod_4906.get(0);
        mod_4905.put(0, t);
    endrule
    rule rule_6330;
        ChannelMessage t;
        t <- mod_4913.get(1);
        mod_4888.put(1, t);
    endrule
    rule rule_6331;
        ChannelMessage t;
        t <- mod_4907.get(1);
        mod_4906.put(1, t);
    endrule
    rule rule_6332;
        ChannelMessage t;
        t <- mod_4892.get(0);
        mod_4893.put(0, t);
    endrule
    rule rule_6333;
        ChannelMessage t;
        t <- mod_4884.get(3);
        mod_4885.put(0, t);
    endrule
    rule rule_6334;
        ChannelMessage t;
        t <- mod_4888.get(0);
        mod_4889.put(0, t);
    endrule
    rule rule_6335;
        ChannelMessage t;
        t <- mod_4891.get(1);
        mod_4892.put(0, t);
    endrule
    rule rule_6336;
        ChannelMessage t;
        t <- mod_4899.get(0);
        mod_4900.put(0, t);
    endrule
    rule rule_6337;
        ChannelMessage t;
        t <- mod_4909.get(0);
        mod_4907.put(0, t);
    endrule
    rule rule_6338;
        ChannelMessage t;
        t <- mod_4886.get(0);
        mod_4911.put(0, t);
    endrule
    rule rule_6339;
        ChannelMessage t;
        t <- mod_4908.get(0);
        mod_4907.put(1, t);
    endrule
    rule rule_6340;
        ChannelMessage t;
        t <- mod_4912.get(0);
        mod_4911.put(1, t);
    endrule
    rule rule_6341;
        ChannelMessage t;
        t <- mod_4911.get(1);
        mod_4906.put(0, t);
    endrule
    rule rule_6342;
        ChannelMessage t;
        t <- mod_4890.get(0);
        mod_4891.put(0, t);
    endrule
    rule rule_6343;
        ChannelMessage t;
        t <- mod_4883.get(1);
        mod_4884.put(0, t);
    endrule
    rule rule_6344;
        ChannelMessage t;
        t <- mod_4882.get(0);
        mod_4883.put(0, t);
    endrule
    rule rule_6345;
        ChannelMessage t;
        t <- mod_4900.get(0);
        mod_4899.put(1, t);
    endrule
    rule rule_6346;
        ChannelMessage t;
        t <- mod_4911.get(0);
        mod_4912.put(0, t);
    endrule
    rule rule_6347;
        ChannelMessage t;
        t <- mod_4887.get(0);
        mod_4917.put(0, t);
    endrule
    rule rule_6348;
        ChannelMessage t;
        t <- mod_4899.get(1);
        mod_4892.put(1, t);
    endrule
    rule rule_6349;
        ChannelMessage t;
        t <- mod_4889.get(0);
        mod_4890.put(0, t);
    endrule
    rule rule_6350;
        ChannelMessage t;
        t <- mod_4904.get(0);
        mod_4890.put(1, t);
    endrule
    rule rule_6351;
        ChannelMessage t;
        t <- mod_4910.get(0);
        mod_4909.put(0, t);
    endrule
    rule rule_6352;
        ChannelMessage t;
        t <- mod_4883.get(0);
        mod_4919.put(0, t);
    endrule
    rule rule_6353;
        ChannelMessage t;
        t <- mod_4898.get(0);
        mod_4898.put(1, t);
    endrule
    rule rule_6354;
        ChannelMessage t;
        t <- mod_4897.get(1);
        mod_4895.put(1, t);
    endrule
    rule rule_6355;
        ChannelMessage t;
        t <- mod_4915.get(0);
        mod_4913.put(0, t);
    endrule
    rule rule_6356;
        ChannelMessage t;
        t <- mod_4895.get(0);
        mod_4897.put(0, t);
    endrule
    rule rule_6357;
        ChannelMessage t;
        t <- mod_4902.get(0);
        mod_4901.put(0, t);
    endrule
    rule rule_6358;
        ChannelMessage t;
        t <- mod_4893.get(0);
        mod_4894.put(0, t);
    endrule
    rule rule_6359;
        ChannelMessage t;
        t <- mod_4881.get(0);
        mod_4882.put(0, t);
    endrule
    rule rule_6360;
        ChannelMessage t;
        t <- mod_4914.get(0);
        mod_4913.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4880.put(0, t);
        end
        if (i == 1) begin
            mod_4896.put(0, t);
        end
        if (i == 2) begin
            mod_4902.put(0, t);
        end
        if (i == 3) begin
            mod_4910.put(0, t);
        end
        if (i == 4) begin
            mod_4916.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_4884.get(0);
        end
        if (i == 2) begin
            t <- mod_4884.get(1);
        end
        if (i == 1) begin
            t <- mod_4884.get(2);
        end
        if (i == 0) begin
            t <- mod_4896.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6154 (Operation_IFC);
    Operation_IFC mod_4921_inner <- mkReshape(2, 64);
    Operation_IFC mod_4921 <- mkDebugOperation(mod_4921_inner, "mod_4921");
    Operation_IFC mod_4922_inner <- mkFlatten(1);
    Operation_IFC mod_4922 <- mkDebugOperation(mod_4922_inner, "mod_4922");
    Operation_IFC mod_4923_inner <- mkFlatten(2);
    Operation_IFC mod_4923 <- mkDebugOperation(mod_4923_inner, "mod_4923");
    Operation_IFC mod_4924_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4924 <- mkDebugOperation(mod_4924_inner, "mod_4924");
    Broadcast_IFC#(4) mod_4925_inner <- mkBroadcast(4);
    Operation_IFC mod_4925 <- mkDebugOperation(mod_4925_inner.op, "mod_4925");
    PMU_IFC mod_4926_bufferize <- mkPMU(2);
    Operation_IFC mod_4926_inner = mod_4926_bufferize.operation;
    Operation_IFC mod_4926 <- mkDebugOperation(mod_4926_inner, "mod_4926");
    Broadcast_IFC#(2) mod_4927_inner <- mkBroadcast(2);
    Operation_IFC mod_4927 <- mkDebugOperation(mod_4927_inner.op, "mod_4927");
    PMU_IFC mod_4928_bufferize <- mkPMU(1);
    Operation_IFC mod_4928_inner = mod_4928_bufferize.operation;
    Operation_IFC mod_4928 <- mkDebugOperation(mod_4928_inner, "mod_4928");
    Operation_IFC mod_4929_inner <- mkBinaryMap(1036, matmul_t_tile);
    Operation_IFC mod_4929 <- mkDebugOperation(mod_4929_inner, "mod_4929");
    Operation_IFC mod_4930_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4930 <- mkDebugOperation(mod_4930_inner, "mod_4930");
    Operation_IFC mod_4931_inner <- mkBinaryMap(1804, mul_tile);
    Operation_IFC mod_4931 <- mkDebugOperation(mod_4931_inner, "mod_4931");
    PMU_IFC mod_4932_bufferize <- mkPMU(1);
    Operation_IFC mod_4932_inner = mod_4932_bufferize.operation;
    Operation_IFC mod_4932 <- mkDebugOperation(mod_4932_inner, "mod_4932");
    Operation_IFC mod_4933_inner <- mkBinaryMap(2323, matmul_t_tile);
    Operation_IFC mod_4933 <- mkDebugOperation(mod_4933_inner, "mod_4933");
    Operation_IFC mod_4934_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4934 <- mkDebugOperation(mod_4934_inner, "mod_4934");
    Operation_IFC mod_4935_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4935 <- mkDebugOperation(mod_4935_inner, "mod_4935");
    Operation_IFC mod_4936_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4936 <- mkDebugOperation(mod_4936_inner, "mod_4936");
    Operation_IFC mod_4937_inner <- mkBinaryMap(2703, mul_tile);
    Operation_IFC mod_4937 <- mkDebugOperation(mod_4937_inner, "mod_4937");
    PMU_IFC mod_4938_bufferize <- mkPMU(1);
    Operation_IFC mod_4938_inner = mod_4938_bufferize.operation;
    Operation_IFC mod_4938 <- mkDebugOperation(mod_4938_inner, "mod_4938");
    PMU_IFC mod_4939_bufferize <- mkPMU(2);
    Operation_IFC mod_4939_inner = mod_4939_bufferize.operation;
    Operation_IFC mod_4939 <- mkDebugOperation(mod_4939_inner, "mod_4939");
    PMU_IFC mod_4940_bufferize <- mkPMU(2);
    Operation_IFC mod_4940_inner = mod_4940_bufferize.operation;
    Operation_IFC mod_4940 <- mkDebugOperation(mod_4940_inner, "mod_4940");
    Operation_IFC mod_4941_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4941 <- mkDebugOperation(mod_4941_inner, "mod_4941");
    Operation_IFC mod_4942_inner <- mkFlatten(1);
    Operation_IFC mod_4942 <- mkDebugOperation(mod_4942_inner, "mod_4942");
    Operation_IFC mod_4943_inner <- mkFlatten(0);
    Operation_IFC mod_4943 <- mkDebugOperation(mod_4943_inner, "mod_4943");
    Operation_IFC mod_4944_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4944 <- mkDebugOperation(mod_4944_inner, "mod_4944");
    Operation_IFC mod_4945_inner <- mkUnaryMap(1676, silu_tile);
    Operation_IFC mod_4945 <- mkDebugOperation(mod_4945_inner, "mod_4945");
    Operation_IFC mod_4946_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4946 <- mkDebugOperation(mod_4946_inner, "mod_4946");
    Operation_IFC mod_4947_inner <- mkBinaryMap(1548, matmul_t_tile);
    Operation_IFC mod_4947 <- mkDebugOperation(mod_4947_inner, "mod_4947");
    PMU_IFC mod_4948_bufferize <- mkPMU(2);
    Operation_IFC mod_4948_inner = mod_4948_bufferize.operation;
    Operation_IFC mod_4948 <- mkDebugOperation(mod_4948_inner, "mod_4948");
    Operation_IFC mod_4949_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4949 <- mkDebugOperation(mod_4949_inner, "mod_4949");
    Operation_IFC mod_4950_inner <- mkFlatten(1);
    Operation_IFC mod_4950 <- mkDebugOperation(mod_4950_inner, "mod_4950");
    Operation_IFC mod_4951_inner <- mkFlatten(0);
    Operation_IFC mod_4951 <- mkDebugOperation(mod_4951_inner, "mod_4951");
    PMU_IFC mod_4952_bufferize <- mkPMU(1);
    Operation_IFC mod_4952_inner = mod_4952_bufferize.operation;
    Operation_IFC mod_4952 <- mkDebugOperation(mod_4952_inner, "mod_4952");
    Operation_IFC mod_4953_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4953 <- mkDebugOperation(mod_4953_inner, "mod_4953");
    PMU_IFC mod_4954_bufferize <- mkPMU(2);
    Operation_IFC mod_4954_inner = mod_4954_bufferize.operation;
    Operation_IFC mod_4954 <- mkDebugOperation(mod_4954_inner, "mod_4954");
    Operation_IFC mod_4955_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4955 <- mkDebugOperation(mod_4955_inner, "mod_4955");
    Operation_IFC mod_4956_inner <- mkFlatten(1);
    Operation_IFC mod_4956 <- mkDebugOperation(mod_4956_inner, "mod_4956");
    Operation_IFC mod_4957_inner <- mkFlatten(0);
    Operation_IFC mod_4957 <- mkDebugOperation(mod_4957_inner, "mod_4957");
    Operation_IFC mod_4958_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4958 <- mkDebugOperation(mod_4958_inner, "mod_4958");
    Operation_IFC mod_4959_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4959 <- mkDebugOperation(mod_4959_inner, "mod_4959");
    PMU_IFC mod_4960_bufferize <- mkPMU(2);
    Operation_IFC mod_4960_inner = mod_4960_bufferize.operation;
    Operation_IFC mod_4960 <- mkDebugOperation(mod_4960_inner, "mod_4960");
    rule rule_6361;
        ChannelMessage t;
        t <- mod_4928.get(1);
        mod_4929.put(0, t);
    endrule
    rule rule_6362;
        ChannelMessage t;
        t <- mod_4929.get(0);
        mod_4930.put(0, t);
    endrule
    rule rule_6363;
        ChannelMessage t;
        t <- mod_4933.get(0);
        mod_4934.put(0, t);
    endrule
    rule rule_6364;
        ChannelMessage t;
        t <- mod_4949.get(0);
        mod_4948.put(1, t);
    endrule
    rule rule_6365;
        ChannelMessage t;
        t <- mod_4958.get(0);
        mod_4928.put(1, t);
    endrule
    rule rule_6366;
        ChannelMessage t;
        t <- mod_4943.get(0);
        mod_4942.put(0, t);
    endrule
    rule rule_6367;
        ChannelMessage t;
        t <- mod_4959.get(0);
        mod_4926.put(1, t);
    endrule
    rule rule_6368;
        ChannelMessage t;
        t <- mod_4940.get(1);
        mod_4933.put(1, t);
    endrule
    rule rule_6369;
        ChannelMessage t;
        t <- mod_4954.get(0);
        mod_4955.put(0, t);
    endrule
    rule rule_6370;
        ChannelMessage t;
        t <- mod_4939.get(0);
        mod_4939.put(1, t);
    endrule
    rule rule_6371;
        ChannelMessage t;
        t <- mod_4946.get(0);
        mod_4945.put(0, t);
    endrule
    rule rule_6372;
        ChannelMessage t;
        t <- mod_4923.get(0);
        mod_4924.put(0, t);
    endrule
    rule rule_6373;
        ChannelMessage t;
        t <- mod_4951.get(0);
        mod_4950.put(0, t);
    endrule
    rule rule_6374;
        ChannelMessage t;
        t <- mod_4952.get(1);
        mod_4947.put(0, t);
    endrule
    rule rule_6375;
        ChannelMessage t;
        t <- mod_4960.get(1);
        mod_4924.put(1, t);
    endrule
    rule rule_6376;
        ChannelMessage t;
        t <- mod_4921.get(0);
        mod_4922.put(0, t);
    endrule
    rule rule_6377;
        ChannelMessage t;
        t <- mod_4924.get(0);
        mod_4960.put(0, t);
    endrule
    rule rule_6378;
        ChannelMessage t;
        t <- mod_4948.get(0);
        mod_4949.put(0, t);
    endrule
    rule rule_6379;
        ChannelMessage t;
        t <- mod_4942.get(0);
        mod_4940.put(0, t);
    endrule
    rule rule_6380;
        ChannelMessage t;
        t <- mod_4928.get(0);
        mod_4958.put(0, t);
    endrule
    rule rule_6381;
        ChannelMessage t;
        t <- mod_4953.get(0);
        mod_4952.put(1, t);
    endrule
    rule rule_6382;
        ChannelMessage t;
        t <- mod_4931.get(0);
        mod_4932.put(0, t);
    endrule
    rule rule_6383;
        ChannelMessage t;
        t <- mod_4941.get(0);
        mod_4940.put(1, t);
    endrule
    rule rule_6384;
        ChannelMessage t;
        t <- mod_4936.get(0);
        mod_4938.put(0, t);
    endrule
    rule rule_6385;
        ChannelMessage t;
        t <- mod_4925.get(3);
        mod_4926.put(0, t);
    endrule
    rule rule_6386;
        ChannelMessage t;
        t <- mod_4927.get(0);
        mod_4952.put(0, t);
    endrule
    rule rule_6387;
        ChannelMessage t;
        t <- mod_4947.get(0);
        mod_4946.put(0, t);
    endrule
    rule rule_6388;
        ChannelMessage t;
        t <- mod_4952.get(0);
        mod_4953.put(0, t);
    endrule
    rule rule_6389;
        ChannelMessage t;
        t <- mod_4954.get(1);
        mod_4929.put(1, t);
    endrule
    rule rule_6390;
        ChannelMessage t;
        t <- mod_4960.get(0);
        mod_4960.put(1, t);
    endrule
    rule rule_6391;
        ChannelMessage t;
        t <- mod_4950.get(0);
        mod_4948.put(0, t);
    endrule
    rule rule_6392;
        ChannelMessage t;
        t <- mod_4922.get(0);
        mod_4923.put(0, t);
    endrule
    rule rule_6393;
        ChannelMessage t;
        t <- mod_4926.get(0);
        mod_4959.put(0, t);
    endrule
    rule rule_6394;
        ChannelMessage t;
        t <- mod_4932.get(0);
        mod_4944.put(0, t);
    endrule
    rule rule_6395;
        ChannelMessage t;
        t <- mod_4936.get(1);
        mod_4937.put(1, t);
    endrule
    rule rule_6396;
        ChannelMessage t;
        t <- mod_4930.get(0);
        mod_4931.put(0, t);
    endrule
    rule rule_6397;
        ChannelMessage t;
        t <- mod_4938.get(1);
        mod_4936.put(1, t);
    endrule
    rule rule_6398;
        ChannelMessage t;
        t <- mod_4932.get(1);
        mod_4933.put(0, t);
    endrule
    rule rule_6399;
        ChannelMessage t;
        t <- mod_4957.get(0);
        mod_4956.put(0, t);
    endrule
    rule rule_6400;
        ChannelMessage t;
        t <- mod_4924.get(1);
        mod_4925.put(0, t);
    endrule
    rule rule_6401;
        ChannelMessage t;
        t <- mod_4935.get(0);
        mod_4939.put(0, t);
    endrule
    rule rule_6402;
        ChannelMessage t;
        t <- mod_4945.get(0);
        mod_4931.put(1, t);
    endrule
    rule rule_6403;
        ChannelMessage t;
        t <- mod_4940.get(0);
        mod_4941.put(0, t);
    endrule
    rule rule_6404;
        ChannelMessage t;
        t <- mod_4927.get(1);
        mod_4928.put(0, t);
    endrule
    rule rule_6405;
        ChannelMessage t;
        t <- mod_4944.get(0);
        mod_4932.put(1, t);
    endrule
    rule rule_6406;
        ChannelMessage t;
        t <- mod_4948.get(1);
        mod_4947.put(1, t);
    endrule
    rule rule_6407;
        ChannelMessage t;
        t <- mod_4934.get(0);
        mod_4935.put(0, t);
    endrule
    rule rule_6408;
        ChannelMessage t;
        t <- mod_4939.get(1);
        mod_4935.put(1, t);
    endrule
    rule rule_6409;
        ChannelMessage t;
        t <- mod_4956.get(0);
        mod_4954.put(0, t);
    endrule
    rule rule_6410;
        ChannelMessage t;
        t <- mod_4926.get(1);
        mod_4927.put(0, t);
    endrule
    rule rule_6411;
        ChannelMessage t;
        t <- mod_4955.get(0);
        mod_4954.put(1, t);
    endrule
    rule rule_6412;
        ChannelMessage t;
        t <- mod_4938.get(0);
        mod_4938.put(1, t);
    endrule
    rule rule_6413;
        ChannelMessage t;
        t <- mod_4935.get(1);
        mod_4936.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4921.put(0, t);
        end
        if (i == 1) begin
            mod_4937.put(0, t);
        end
        if (i == 2) begin
            mod_4943.put(0, t);
        end
        if (i == 3) begin
            mod_4951.put(0, t);
        end
        if (i == 4) begin
            mod_4957.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 2) begin
            t <- mod_4925.get(0);
        end
        if (i == 1) begin
            t <- mod_4925.get(1);
        end
        if (i == 0) begin
            t <- mod_4925.get(2);
        end
        if (i == 3) begin
            t <- mod_4937.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6155 (Operation_IFC);
    Operation_IFC mod_4962_inner <- mkReshape(2, 64);
    Operation_IFC mod_4962 <- mkDebugOperation(mod_4962_inner, "mod_4962");
    Operation_IFC mod_4963_inner <- mkFlatten(1);
    Operation_IFC mod_4963 <- mkDebugOperation(mod_4963_inner, "mod_4963");
    Operation_IFC mod_4964_inner <- mkFlatten(2);
    Operation_IFC mod_4964 <- mkDebugOperation(mod_4964_inner, "mod_4964");
    Operation_IFC mod_4965_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4965 <- mkDebugOperation(mod_4965_inner, "mod_4965");
    Broadcast_IFC#(4) mod_4966_inner <- mkBroadcast(4);
    Operation_IFC mod_4966 <- mkDebugOperation(mod_4966_inner.op, "mod_4966");
    PMU_IFC mod_4967_bufferize <- mkPMU(2);
    Operation_IFC mod_4967_inner = mod_4967_bufferize.operation;
    Operation_IFC mod_4967 <- mkDebugOperation(mod_4967_inner, "mod_4967");
    Broadcast_IFC#(2) mod_4968_inner <- mkBroadcast(2);
    Operation_IFC mod_4968 <- mkDebugOperation(mod_4968_inner.op, "mod_4968");
    PMU_IFC mod_4969_bufferize <- mkPMU(1);
    Operation_IFC mod_4969_inner = mod_4969_bufferize.operation;
    Operation_IFC mod_4969 <- mkDebugOperation(mod_4969_inner, "mod_4969");
    Operation_IFC mod_4970_inner <- mkBinaryMap(1035, matmul_t_tile);
    Operation_IFC mod_4970 <- mkDebugOperation(mod_4970_inner, "mod_4970");
    Operation_IFC mod_4971_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4971 <- mkDebugOperation(mod_4971_inner, "mod_4971");
    Operation_IFC mod_4972_inner <- mkBinaryMap(1803, mul_tile);
    Operation_IFC mod_4972 <- mkDebugOperation(mod_4972_inner, "mod_4972");
    PMU_IFC mod_4973_bufferize <- mkPMU(1);
    Operation_IFC mod_4973_inner = mod_4973_bufferize.operation;
    Operation_IFC mod_4973 <- mkDebugOperation(mod_4973_inner, "mod_4973");
    Operation_IFC mod_4974_inner <- mkBinaryMap(2321, matmul_t_tile);
    Operation_IFC mod_4974 <- mkDebugOperation(mod_4974_inner, "mod_4974");
    Operation_IFC mod_4975_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4975 <- mkDebugOperation(mod_4975_inner, "mod_4975");
    Operation_IFC mod_4976_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4976 <- mkDebugOperation(mod_4976_inner, "mod_4976");
    Operation_IFC mod_4977_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4977 <- mkDebugOperation(mod_4977_inner, "mod_4977");
    Operation_IFC mod_4978_inner <- mkBinaryMap(2702, mul_tile);
    Operation_IFC mod_4978 <- mkDebugOperation(mod_4978_inner, "mod_4978");
    PMU_IFC mod_4979_bufferize <- mkPMU(1);
    Operation_IFC mod_4979_inner = mod_4979_bufferize.operation;
    Operation_IFC mod_4979 <- mkDebugOperation(mod_4979_inner, "mod_4979");
    PMU_IFC mod_4980_bufferize <- mkPMU(2);
    Operation_IFC mod_4980_inner = mod_4980_bufferize.operation;
    Operation_IFC mod_4980 <- mkDebugOperation(mod_4980_inner, "mod_4980");
    PMU_IFC mod_4981_bufferize <- mkPMU(2);
    Operation_IFC mod_4981_inner = mod_4981_bufferize.operation;
    Operation_IFC mod_4981 <- mkDebugOperation(mod_4981_inner, "mod_4981");
    Operation_IFC mod_4982_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4982 <- mkDebugOperation(mod_4982_inner, "mod_4982");
    Operation_IFC mod_4983_inner <- mkFlatten(1);
    Operation_IFC mod_4983 <- mkDebugOperation(mod_4983_inner, "mod_4983");
    Operation_IFC mod_4984_inner <- mkFlatten(0);
    Operation_IFC mod_4984 <- mkDebugOperation(mod_4984_inner, "mod_4984");
    Operation_IFC mod_4985_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4985 <- mkDebugOperation(mod_4985_inner, "mod_4985");
    Operation_IFC mod_4986_inner <- mkUnaryMap(1675, silu_tile);
    Operation_IFC mod_4986 <- mkDebugOperation(mod_4986_inner, "mod_4986");
    Operation_IFC mod_4987_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4987 <- mkDebugOperation(mod_4987_inner, "mod_4987");
    Operation_IFC mod_4988_inner <- mkBinaryMap(1547, matmul_t_tile);
    Operation_IFC mod_4988 <- mkDebugOperation(mod_4988_inner, "mod_4988");
    PMU_IFC mod_4989_bufferize <- mkPMU(2);
    Operation_IFC mod_4989_inner = mod_4989_bufferize.operation;
    Operation_IFC mod_4989 <- mkDebugOperation(mod_4989_inner, "mod_4989");
    Operation_IFC mod_4990_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4990 <- mkDebugOperation(mod_4990_inner, "mod_4990");
    Operation_IFC mod_4991_inner <- mkFlatten(1);
    Operation_IFC mod_4991 <- mkDebugOperation(mod_4991_inner, "mod_4991");
    Operation_IFC mod_4992_inner <- mkFlatten(0);
    Operation_IFC mod_4992 <- mkDebugOperation(mod_4992_inner, "mod_4992");
    PMU_IFC mod_4993_bufferize <- mkPMU(1);
    Operation_IFC mod_4993_inner = mod_4993_bufferize.operation;
    Operation_IFC mod_4993 <- mkDebugOperation(mod_4993_inner, "mod_4993");
    Operation_IFC mod_4994_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4994 <- mkDebugOperation(mod_4994_inner, "mod_4994");
    PMU_IFC mod_4995_bufferize <- mkPMU(2);
    Operation_IFC mod_4995_inner = mod_4995_bufferize.operation;
    Operation_IFC mod_4995 <- mkDebugOperation(mod_4995_inner, "mod_4995");
    Operation_IFC mod_4996_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4996 <- mkDebugOperation(mod_4996_inner, "mod_4996");
    Operation_IFC mod_4997_inner <- mkFlatten(1);
    Operation_IFC mod_4997 <- mkDebugOperation(mod_4997_inner, "mod_4997");
    Operation_IFC mod_4998_inner <- mkFlatten(0);
    Operation_IFC mod_4998 <- mkDebugOperation(mod_4998_inner, "mod_4998");
    Operation_IFC mod_4999_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4999 <- mkDebugOperation(mod_4999_inner, "mod_4999");
    Operation_IFC mod_5000_inner <- mkRepeatStatic(2);
    Operation_IFC mod_5000 <- mkDebugOperation(mod_5000_inner, "mod_5000");
    PMU_IFC mod_5001_bufferize <- mkPMU(2);
    Operation_IFC mod_5001_inner = mod_5001_bufferize.operation;
    Operation_IFC mod_5001 <- mkDebugOperation(mod_5001_inner, "mod_5001");
    rule rule_6414;
        ChannelMessage t;
        t <- mod_4962.get(0);
        mod_4963.put(0, t);
    endrule
    rule rule_6415;
        ChannelMessage t;
        t <- mod_4979.get(0);
        mod_4979.put(1, t);
    endrule
    rule rule_6416;
        ChannelMessage t;
        t <- mod_4993.get(0);
        mod_4994.put(0, t);
    endrule
    rule rule_6417;
        ChannelMessage t;
        t <- mod_5001.get(0);
        mod_5001.put(1, t);
    endrule
    rule rule_6418;
        ChannelMessage t;
        t <- mod_4973.get(0);
        mod_4985.put(0, t);
    endrule
    rule rule_6419;
        ChannelMessage t;
        t <- mod_4998.get(0);
        mod_4997.put(0, t);
    endrule
    rule rule_6420;
        ChannelMessage t;
        t <- mod_4999.get(0);
        mod_4969.put(1, t);
    endrule
    rule rule_6421;
        ChannelMessage t;
        t <- mod_4995.get(0);
        mod_4996.put(0, t);
    endrule
    rule rule_6422;
        ChannelMessage t;
        t <- mod_4968.get(0);
        mod_4993.put(0, t);
    endrule
    rule rule_6423;
        ChannelMessage t;
        t <- mod_4969.get(0);
        mod_4999.put(0, t);
    endrule
    rule rule_6424;
        ChannelMessage t;
        t <- mod_4968.get(1);
        mod_4969.put(0, t);
    endrule
    rule rule_6425;
        ChannelMessage t;
        t <- mod_4989.get(1);
        mod_4988.put(1, t);
    endrule
    rule rule_6426;
        ChannelMessage t;
        t <- mod_4980.get(0);
        mod_4980.put(1, t);
    endrule
    rule rule_6427;
        ChannelMessage t;
        t <- mod_4985.get(0);
        mod_4973.put(1, t);
    endrule
    rule rule_6428;
        ChannelMessage t;
        t <- mod_4970.get(0);
        mod_4971.put(0, t);
    endrule
    rule rule_6429;
        ChannelMessage t;
        t <- mod_5000.get(0);
        mod_4967.put(1, t);
    endrule
    rule rule_6430;
        ChannelMessage t;
        t <- mod_4991.get(0);
        mod_4989.put(0, t);
    endrule
    rule rule_6431;
        ChannelMessage t;
        t <- mod_4988.get(0);
        mod_4987.put(0, t);
    endrule
    rule rule_6432;
        ChannelMessage t;
        t <- mod_4983.get(0);
        mod_4981.put(0, t);
    endrule
    rule rule_6433;
        ChannelMessage t;
        t <- mod_4997.get(0);
        mod_4995.put(0, t);
    endrule
    rule rule_6434;
        ChannelMessage t;
        t <- mod_4976.get(1);
        mod_4977.put(0, t);
    endrule
    rule rule_6435;
        ChannelMessage t;
        t <- mod_4981.get(0);
        mod_4982.put(0, t);
    endrule
    rule rule_6436;
        ChannelMessage t;
        t <- mod_4969.get(1);
        mod_4970.put(0, t);
    endrule
    rule rule_6437;
        ChannelMessage t;
        t <- mod_4974.get(0);
        mod_4975.put(0, t);
    endrule
    rule rule_6438;
        ChannelMessage t;
        t <- mod_4993.get(1);
        mod_4988.put(0, t);
    endrule
    rule rule_6439;
        ChannelMessage t;
        t <- mod_4982.get(0);
        mod_4981.put(1, t);
    endrule
    rule rule_6440;
        ChannelMessage t;
        t <- mod_4971.get(0);
        mod_4972.put(0, t);
    endrule
    rule rule_6441;
        ChannelMessage t;
        t <- mod_4967.get(1);
        mod_4968.put(0, t);
    endrule
    rule rule_6442;
        ChannelMessage t;
        t <- mod_4972.get(0);
        mod_4973.put(0, t);
    endrule
    rule rule_6443;
        ChannelMessage t;
        t <- mod_4981.get(1);
        mod_4974.put(1, t);
    endrule
    rule rule_6444;
        ChannelMessage t;
        t <- mod_4965.get(0);
        mod_5001.put(0, t);
    endrule
    rule rule_6445;
        ChannelMessage t;
        t <- mod_4976.get(0);
        mod_4980.put(0, t);
    endrule
    rule rule_6446;
        ChannelMessage t;
        t <- mod_4984.get(0);
        mod_4983.put(0, t);
    endrule
    rule rule_6447;
        ChannelMessage t;
        t <- mod_4965.get(1);
        mod_4966.put(0, t);
    endrule
    rule rule_6448;
        ChannelMessage t;
        t <- mod_4977.get(1);
        mod_4978.put(1, t);
    endrule
    rule rule_6449;
        ChannelMessage t;
        t <- mod_4986.get(0);
        mod_4972.put(1, t);
    endrule
    rule rule_6450;
        ChannelMessage t;
        t <- mod_4994.get(0);
        mod_4993.put(1, t);
    endrule
    rule rule_6451;
        ChannelMessage t;
        t <- mod_4989.get(0);
        mod_4990.put(0, t);
    endrule
    rule rule_6452;
        ChannelMessage t;
        t <- mod_4964.get(0);
        mod_4965.put(0, t);
    endrule
    rule rule_6453;
        ChannelMessage t;
        t <- mod_4979.get(1);
        mod_4977.put(1, t);
    endrule
    rule rule_6454;
        ChannelMessage t;
        t <- mod_4963.get(0);
        mod_4964.put(0, t);
    endrule
    rule rule_6455;
        ChannelMessage t;
        t <- mod_4967.get(0);
        mod_5000.put(0, t);
    endrule
    rule rule_6456;
        ChannelMessage t;
        t <- mod_4973.get(1);
        mod_4974.put(0, t);
    endrule
    rule rule_6457;
        ChannelMessage t;
        t <- mod_4975.get(0);
        mod_4976.put(0, t);
    endrule
    rule rule_6458;
        ChannelMessage t;
        t <- mod_4977.get(0);
        mod_4979.put(0, t);
    endrule
    rule rule_6459;
        ChannelMessage t;
        t <- mod_4996.get(0);
        mod_4995.put(1, t);
    endrule
    rule rule_6460;
        ChannelMessage t;
        t <- mod_4990.get(0);
        mod_4989.put(1, t);
    endrule
    rule rule_6461;
        ChannelMessage t;
        t <- mod_4987.get(0);
        mod_4986.put(0, t);
    endrule
    rule rule_6462;
        ChannelMessage t;
        t <- mod_4992.get(0);
        mod_4991.put(0, t);
    endrule
    rule rule_6463;
        ChannelMessage t;
        t <- mod_4966.get(3);
        mod_4967.put(0, t);
    endrule
    rule rule_6464;
        ChannelMessage t;
        t <- mod_4995.get(1);
        mod_4970.put(1, t);
    endrule
    rule rule_6465;
        ChannelMessage t;
        t <- mod_5001.get(1);
        mod_4965.put(1, t);
    endrule
    rule rule_6466;
        ChannelMessage t;
        t <- mod_4980.get(1);
        mod_4976.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4962.put(0, t);
        end
        if (i == 1) begin
            mod_4978.put(0, t);
        end
        if (i == 2) begin
            mod_4984.put(0, t);
        end
        if (i == 3) begin
            mod_4992.put(0, t);
        end
        if (i == 4) begin
            mod_4998.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_4966.get(0);
        end
        if (i == 1) begin
            t <- mod_4966.get(1);
        end
        if (i == 0) begin
            t <- mod_4966.get(2);
        end
        if (i == 2) begin
            t <- mod_4978.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6156 (Operation_IFC);
    Operation_IFC mod_5003_inner <- mkReshape(2, 64);
    Operation_IFC mod_5003 <- mkDebugOperation(mod_5003_inner, "mod_5003");
    Operation_IFC mod_5004_inner <- mkFlatten(1);
    Operation_IFC mod_5004 <- mkDebugOperation(mod_5004_inner, "mod_5004");
    Operation_IFC mod_5005_inner <- mkFlatten(2);
    Operation_IFC mod_5005 <- mkDebugOperation(mod_5005_inner, "mod_5005");
    Operation_IFC mod_5006_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_5006 <- mkDebugOperation(mod_5006_inner, "mod_5006");
    Broadcast_IFC#(4) mod_5007_inner <- mkBroadcast(4);
    Operation_IFC mod_5007 <- mkDebugOperation(mod_5007_inner.op, "mod_5007");
    PMU_IFC mod_5008_bufferize <- mkPMU(2);
    Operation_IFC mod_5008_inner = mod_5008_bufferize.operation;
    Operation_IFC mod_5008 <- mkDebugOperation(mod_5008_inner, "mod_5008");
    Broadcast_IFC#(2) mod_5009_inner <- mkBroadcast(2);
    Operation_IFC mod_5009 <- mkDebugOperation(mod_5009_inner.op, "mod_5009");
    PMU_IFC mod_5010_bufferize <- mkPMU(1);
    Operation_IFC mod_5010_inner = mod_5010_bufferize.operation;
    Operation_IFC mod_5010 <- mkDebugOperation(mod_5010_inner, "mod_5010");
    Operation_IFC mod_5011_inner <- mkBinaryMap(1034, matmul_t_tile);
    Operation_IFC mod_5011 <- mkDebugOperation(mod_5011_inner, "mod_5011");
    Operation_IFC mod_5012_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_5012 <- mkDebugOperation(mod_5012_inner, "mod_5012");
    Operation_IFC mod_5013_inner <- mkBinaryMap(1802, mul_tile);
    Operation_IFC mod_5013 <- mkDebugOperation(mod_5013_inner, "mod_5013");
    PMU_IFC mod_5014_bufferize <- mkPMU(1);
    Operation_IFC mod_5014_inner = mod_5014_bufferize.operation;
    Operation_IFC mod_5014 <- mkDebugOperation(mod_5014_inner, "mod_5014");
    Operation_IFC mod_5015_inner <- mkBinaryMap(2319, matmul_t_tile);
    Operation_IFC mod_5015 <- mkDebugOperation(mod_5015_inner, "mod_5015");
    Operation_IFC mod_5016_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_5016 <- mkDebugOperation(mod_5016_inner, "mod_5016");
    Operation_IFC mod_5017_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_5017 <- mkDebugOperation(mod_5017_inner, "mod_5017");
    Operation_IFC mod_5018_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_5018 <- mkDebugOperation(mod_5018_inner, "mod_5018");
    Operation_IFC mod_5019_inner <- mkBinaryMap(2701, mul_tile);
    Operation_IFC mod_5019 <- mkDebugOperation(mod_5019_inner, "mod_5019");
    PMU_IFC mod_5020_bufferize <- mkPMU(1);
    Operation_IFC mod_5020_inner = mod_5020_bufferize.operation;
    Operation_IFC mod_5020 <- mkDebugOperation(mod_5020_inner, "mod_5020");
    PMU_IFC mod_5021_bufferize <- mkPMU(2);
    Operation_IFC mod_5021_inner = mod_5021_bufferize.operation;
    Operation_IFC mod_5021 <- mkDebugOperation(mod_5021_inner, "mod_5021");
    PMU_IFC mod_5022_bufferize <- mkPMU(2);
    Operation_IFC mod_5022_inner = mod_5022_bufferize.operation;
    Operation_IFC mod_5022 <- mkDebugOperation(mod_5022_inner, "mod_5022");
    Operation_IFC mod_5023_inner <- mkRepeatStatic(8);
    Operation_IFC mod_5023 <- mkDebugOperation(mod_5023_inner, "mod_5023");
    Operation_IFC mod_5024_inner <- mkFlatten(1);
    Operation_IFC mod_5024 <- mkDebugOperation(mod_5024_inner, "mod_5024");
    Operation_IFC mod_5025_inner <- mkFlatten(0);
    Operation_IFC mod_5025 <- mkDebugOperation(mod_5025_inner, "mod_5025");
    Operation_IFC mod_5026_inner <- mkRepeatStatic(3);
    Operation_IFC mod_5026 <- mkDebugOperation(mod_5026_inner, "mod_5026");
    Operation_IFC mod_5027_inner <- mkUnaryMap(1674, silu_tile);
    Operation_IFC mod_5027 <- mkDebugOperation(mod_5027_inner, "mod_5027");
    Operation_IFC mod_5028_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_5028 <- mkDebugOperation(mod_5028_inner, "mod_5028");
    Operation_IFC mod_5029_inner <- mkBinaryMap(1546, matmul_t_tile);
    Operation_IFC mod_5029 <- mkDebugOperation(mod_5029_inner, "mod_5029");
    PMU_IFC mod_5030_bufferize <- mkPMU(2);
    Operation_IFC mod_5030_inner = mod_5030_bufferize.operation;
    Operation_IFC mod_5030 <- mkDebugOperation(mod_5030_inner, "mod_5030");
    Operation_IFC mod_5031_inner <- mkRepeatStatic(8);
    Operation_IFC mod_5031 <- mkDebugOperation(mod_5031_inner, "mod_5031");
    Operation_IFC mod_5032_inner <- mkFlatten(1);
    Operation_IFC mod_5032 <- mkDebugOperation(mod_5032_inner, "mod_5032");
    Operation_IFC mod_5033_inner <- mkFlatten(0);
    Operation_IFC mod_5033 <- mkDebugOperation(mod_5033_inner, "mod_5033");
    PMU_IFC mod_5034_bufferize <- mkPMU(1);
    Operation_IFC mod_5034_inner = mod_5034_bufferize.operation;
    Operation_IFC mod_5034 <- mkDebugOperation(mod_5034_inner, "mod_5034");
    Operation_IFC mod_5035_inner <- mkRepeatStatic(16);
    Operation_IFC mod_5035 <- mkDebugOperation(mod_5035_inner, "mod_5035");
    PMU_IFC mod_5036_bufferize <- mkPMU(2);
    Operation_IFC mod_5036_inner = mod_5036_bufferize.operation;
    Operation_IFC mod_5036 <- mkDebugOperation(mod_5036_inner, "mod_5036");
    Operation_IFC mod_5037_inner <- mkRepeatStatic(8);
    Operation_IFC mod_5037 <- mkDebugOperation(mod_5037_inner, "mod_5037");
    Operation_IFC mod_5038_inner <- mkFlatten(1);
    Operation_IFC mod_5038 <- mkDebugOperation(mod_5038_inner, "mod_5038");
    Operation_IFC mod_5039_inner <- mkFlatten(0);
    Operation_IFC mod_5039 <- mkDebugOperation(mod_5039_inner, "mod_5039");
    Operation_IFC mod_5040_inner <- mkRepeatStatic(16);
    Operation_IFC mod_5040 <- mkDebugOperation(mod_5040_inner, "mod_5040");
    Operation_IFC mod_5041_inner <- mkRepeatStatic(2);
    Operation_IFC mod_5041 <- mkDebugOperation(mod_5041_inner, "mod_5041");
    PMU_IFC mod_5042_bufferize <- mkPMU(2);
    Operation_IFC mod_5042_inner = mod_5042_bufferize.operation;
    Operation_IFC mod_5042 <- mkDebugOperation(mod_5042_inner, "mod_5042");
    rule rule_6467;
        ChannelMessage t;
        t <- mod_5006.get(1);
        mod_5007.put(0, t);
    endrule
    rule rule_6468;
        ChannelMessage t;
        t <- mod_5029.get(0);
        mod_5028.put(0, t);
    endrule
    rule rule_6469;
        ChannelMessage t;
        t <- mod_5020.get(1);
        mod_5018.put(1, t);
    endrule
    rule rule_6470;
        ChannelMessage t;
        t <- mod_5022.get(0);
        mod_5023.put(0, t);
    endrule
    rule rule_6471;
        ChannelMessage t;
        t <- mod_5032.get(0);
        mod_5030.put(0, t);
    endrule
    rule rule_6472;
        ChannelMessage t;
        t <- mod_5017.get(0);
        mod_5021.put(0, t);
    endrule
    rule rule_6473;
        ChannelMessage t;
        t <- mod_5007.get(3);
        mod_5008.put(0, t);
    endrule
    rule rule_6474;
        ChannelMessage t;
        t <- mod_5021.get(1);
        mod_5017.put(1, t);
    endrule
    rule rule_6475;
        ChannelMessage t;
        t <- mod_5024.get(0);
        mod_5022.put(0, t);
    endrule
    rule rule_6476;
        ChannelMessage t;
        t <- mod_5037.get(0);
        mod_5036.put(1, t);
    endrule
    rule rule_6477;
        ChannelMessage t;
        t <- mod_5022.get(1);
        mod_5015.put(1, t);
    endrule
    rule rule_6478;
        ChannelMessage t;
        t <- mod_5027.get(0);
        mod_5013.put(1, t);
    endrule
    rule rule_6479;
        ChannelMessage t;
        t <- mod_5042.get(0);
        mod_5042.put(1, t);
    endrule
    rule rule_6480;
        ChannelMessage t;
        t <- mod_5017.get(1);
        mod_5018.put(0, t);
    endrule
    rule rule_6481;
        ChannelMessage t;
        t <- mod_5025.get(0);
        mod_5024.put(0, t);
    endrule
    rule rule_6482;
        ChannelMessage t;
        t <- mod_5016.get(0);
        mod_5017.put(0, t);
    endrule
    rule rule_6483;
        ChannelMessage t;
        t <- mod_5026.get(0);
        mod_5014.put(1, t);
    endrule
    rule rule_6484;
        ChannelMessage t;
        t <- mod_5010.get(0);
        mod_5040.put(0, t);
    endrule
    rule rule_6485;
        ChannelMessage t;
        t <- mod_5011.get(0);
        mod_5012.put(0, t);
    endrule
    rule rule_6486;
        ChannelMessage t;
        t <- mod_5013.get(0);
        mod_5014.put(0, t);
    endrule
    rule rule_6487;
        ChannelMessage t;
        t <- mod_5003.get(0);
        mod_5004.put(0, t);
    endrule
    rule rule_6488;
        ChannelMessage t;
        t <- mod_5006.get(0);
        mod_5042.put(0, t);
    endrule
    rule rule_6489;
        ChannelMessage t;
        t <- mod_5042.get(1);
        mod_5006.put(1, t);
    endrule
    rule rule_6490;
        ChannelMessage t;
        t <- mod_5035.get(0);
        mod_5034.put(1, t);
    endrule
    rule rule_6491;
        ChannelMessage t;
        t <- mod_5028.get(0);
        mod_5027.put(0, t);
    endrule
    rule rule_6492;
        ChannelMessage t;
        t <- mod_5014.get(0);
        mod_5026.put(0, t);
    endrule
    rule rule_6493;
        ChannelMessage t;
        t <- mod_5030.get(1);
        mod_5029.put(1, t);
    endrule
    rule rule_6494;
        ChannelMessage t;
        t <- mod_5012.get(0);
        mod_5013.put(0, t);
    endrule
    rule rule_6495;
        ChannelMessage t;
        t <- mod_5021.get(0);
        mod_5021.put(1, t);
    endrule
    rule rule_6496;
        ChannelMessage t;
        t <- mod_5038.get(0);
        mod_5036.put(0, t);
    endrule
    rule rule_6497;
        ChannelMessage t;
        t <- mod_5008.get(0);
        mod_5041.put(0, t);
    endrule
    rule rule_6498;
        ChannelMessage t;
        t <- mod_5008.get(1);
        mod_5009.put(0, t);
    endrule
    rule rule_6499;
        ChannelMessage t;
        t <- mod_5004.get(0);
        mod_5005.put(0, t);
    endrule
    rule rule_6500;
        ChannelMessage t;
        t <- mod_5010.get(1);
        mod_5011.put(0, t);
    endrule
    rule rule_6501;
        ChannelMessage t;
        t <- mod_5018.get(1);
        mod_5019.put(1, t);
    endrule
    rule rule_6502;
        ChannelMessage t;
        t <- mod_5023.get(0);
        mod_5022.put(1, t);
    endrule
    rule rule_6503;
        ChannelMessage t;
        t <- mod_5015.get(0);
        mod_5016.put(0, t);
    endrule
    rule rule_6504;
        ChannelMessage t;
        t <- mod_5034.get(1);
        mod_5029.put(0, t);
    endrule
    rule rule_6505;
        ChannelMessage t;
        t <- mod_5039.get(0);
        mod_5038.put(0, t);
    endrule
    rule rule_6506;
        ChannelMessage t;
        t <- mod_5036.get(0);
        mod_5037.put(0, t);
    endrule
    rule rule_6507;
        ChannelMessage t;
        t <- mod_5009.get(1);
        mod_5010.put(0, t);
    endrule
    rule rule_6508;
        ChannelMessage t;
        t <- mod_5014.get(1);
        mod_5015.put(0, t);
    endrule
    rule rule_6509;
        ChannelMessage t;
        t <- mod_5034.get(0);
        mod_5035.put(0, t);
    endrule
    rule rule_6510;
        ChannelMessage t;
        t <- mod_5036.get(1);
        mod_5011.put(1, t);
    endrule
    rule rule_6511;
        ChannelMessage t;
        t <- mod_5031.get(0);
        mod_5030.put(1, t);
    endrule
    rule rule_6512;
        ChannelMessage t;
        t <- mod_5033.get(0);
        mod_5032.put(0, t);
    endrule
    rule rule_6513;
        ChannelMessage t;
        t <- mod_5040.get(0);
        mod_5010.put(1, t);
    endrule
    rule rule_6514;
        ChannelMessage t;
        t <- mod_5041.get(0);
        mod_5008.put(1, t);
    endrule
    rule rule_6515;
        ChannelMessage t;
        t <- mod_5018.get(0);
        mod_5020.put(0, t);
    endrule
    rule rule_6516;
        ChannelMessage t;
        t <- mod_5005.get(0);
        mod_5006.put(0, t);
    endrule
    rule rule_6517;
        ChannelMessage t;
        t <- mod_5020.get(0);
        mod_5020.put(1, t);
    endrule
    rule rule_6518;
        ChannelMessage t;
        t <- mod_5030.get(0);
        mod_5031.put(0, t);
    endrule
    rule rule_6519;
        ChannelMessage t;
        t <- mod_5009.get(0);
        mod_5034.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_5003.put(0, t);
        end
        if (i == 1) begin
            mod_5019.put(0, t);
        end
        if (i == 2) begin
            mod_5025.put(0, t);
        end
        if (i == 3) begin
            mod_5033.put(0, t);
        end
        if (i == 4) begin
            mod_5039.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_5007.get(0);
        end
        if (i == 2) begin
            t <- mod_5007.get(1);
        end
        if (i == 3) begin
            t <- mod_5007.get(2);
        end
        if (i == 0) begin
            t <- mod_5019.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6157 (Operation_IFC);
    Operation_IFC mod_5044_inner <- mkReshape(2, 64);
    Operation_IFC mod_5044 <- mkDebugOperation(mod_5044_inner, "mod_5044");
    Operation_IFC mod_5045_inner <- mkFlatten(1);
    Operation_IFC mod_5045 <- mkDebugOperation(mod_5045_inner, "mod_5045");
    Operation_IFC mod_5046_inner <- mkFlatten(2);
    Operation_IFC mod_5046 <- mkDebugOperation(mod_5046_inner, "mod_5046");
    Operation_IFC mod_5047_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_5047 <- mkDebugOperation(mod_5047_inner, "mod_5047");
    Broadcast_IFC#(4) mod_5048_inner <- mkBroadcast(4);
    Operation_IFC mod_5048 <- mkDebugOperation(mod_5048_inner.op, "mod_5048");
    PMU_IFC mod_5049_bufferize <- mkPMU(2);
    Operation_IFC mod_5049_inner = mod_5049_bufferize.operation;
    Operation_IFC mod_5049 <- mkDebugOperation(mod_5049_inner, "mod_5049");
    Broadcast_IFC#(2) mod_5050_inner <- mkBroadcast(2);
    Operation_IFC mod_5050 <- mkDebugOperation(mod_5050_inner.op, "mod_5050");
    PMU_IFC mod_5051_bufferize <- mkPMU(1);
    Operation_IFC mod_5051_inner = mod_5051_bufferize.operation;
    Operation_IFC mod_5051 <- mkDebugOperation(mod_5051_inner, "mod_5051");
    Operation_IFC mod_5052_inner <- mkBinaryMap(1033, matmul_t_tile);
    Operation_IFC mod_5052 <- mkDebugOperation(mod_5052_inner, "mod_5052");
    Operation_IFC mod_5053_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_5053 <- mkDebugOperation(mod_5053_inner, "mod_5053");
    Operation_IFC mod_5054_inner <- mkBinaryMap(1801, mul_tile);
    Operation_IFC mod_5054 <- mkDebugOperation(mod_5054_inner, "mod_5054");
    PMU_IFC mod_5055_bufferize <- mkPMU(1);
    Operation_IFC mod_5055_inner = mod_5055_bufferize.operation;
    Operation_IFC mod_5055 <- mkDebugOperation(mod_5055_inner, "mod_5055");
    Operation_IFC mod_5056_inner <- mkBinaryMap(2317, matmul_t_tile);
    Operation_IFC mod_5056 <- mkDebugOperation(mod_5056_inner, "mod_5056");
    Operation_IFC mod_5057_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_5057 <- mkDebugOperation(mod_5057_inner, "mod_5057");
    Operation_IFC mod_5058_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_5058 <- mkDebugOperation(mod_5058_inner, "mod_5058");
    Operation_IFC mod_5059_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_5059 <- mkDebugOperation(mod_5059_inner, "mod_5059");
    Operation_IFC mod_5060_inner <- mkBinaryMap(2700, mul_tile);
    Operation_IFC mod_5060 <- mkDebugOperation(mod_5060_inner, "mod_5060");
    PMU_IFC mod_5061_bufferize <- mkPMU(1);
    Operation_IFC mod_5061_inner = mod_5061_bufferize.operation;
    Operation_IFC mod_5061 <- mkDebugOperation(mod_5061_inner, "mod_5061");
    PMU_IFC mod_5062_bufferize <- mkPMU(2);
    Operation_IFC mod_5062_inner = mod_5062_bufferize.operation;
    Operation_IFC mod_5062 <- mkDebugOperation(mod_5062_inner, "mod_5062");
    PMU_IFC mod_5063_bufferize <- mkPMU(2);
    Operation_IFC mod_5063_inner = mod_5063_bufferize.operation;
    Operation_IFC mod_5063 <- mkDebugOperation(mod_5063_inner, "mod_5063");
    Operation_IFC mod_5064_inner <- mkRepeatStatic(8);
    Operation_IFC mod_5064 <- mkDebugOperation(mod_5064_inner, "mod_5064");
    Operation_IFC mod_5065_inner <- mkFlatten(1);
    Operation_IFC mod_5065 <- mkDebugOperation(mod_5065_inner, "mod_5065");
    Operation_IFC mod_5066_inner <- mkFlatten(0);
    Operation_IFC mod_5066 <- mkDebugOperation(mod_5066_inner, "mod_5066");
    Operation_IFC mod_5067_inner <- mkRepeatStatic(3);
    Operation_IFC mod_5067 <- mkDebugOperation(mod_5067_inner, "mod_5067");
    Operation_IFC mod_5068_inner <- mkUnaryMap(1673, silu_tile);
    Operation_IFC mod_5068 <- mkDebugOperation(mod_5068_inner, "mod_5068");
    Operation_IFC mod_5069_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_5069 <- mkDebugOperation(mod_5069_inner, "mod_5069");
    Operation_IFC mod_5070_inner <- mkBinaryMap(1545, matmul_t_tile);
    Operation_IFC mod_5070 <- mkDebugOperation(mod_5070_inner, "mod_5070");
    PMU_IFC mod_5071_bufferize <- mkPMU(2);
    Operation_IFC mod_5071_inner = mod_5071_bufferize.operation;
    Operation_IFC mod_5071 <- mkDebugOperation(mod_5071_inner, "mod_5071");
    Operation_IFC mod_5072_inner <- mkRepeatStatic(8);
    Operation_IFC mod_5072 <- mkDebugOperation(mod_5072_inner, "mod_5072");
    Operation_IFC mod_5073_inner <- mkFlatten(1);
    Operation_IFC mod_5073 <- mkDebugOperation(mod_5073_inner, "mod_5073");
    Operation_IFC mod_5074_inner <- mkFlatten(0);
    Operation_IFC mod_5074 <- mkDebugOperation(mod_5074_inner, "mod_5074");
    PMU_IFC mod_5075_bufferize <- mkPMU(1);
    Operation_IFC mod_5075_inner = mod_5075_bufferize.operation;
    Operation_IFC mod_5075 <- mkDebugOperation(mod_5075_inner, "mod_5075");
    Operation_IFC mod_5076_inner <- mkRepeatStatic(16);
    Operation_IFC mod_5076 <- mkDebugOperation(mod_5076_inner, "mod_5076");
    PMU_IFC mod_5077_bufferize <- mkPMU(2);
    Operation_IFC mod_5077_inner = mod_5077_bufferize.operation;
    Operation_IFC mod_5077 <- mkDebugOperation(mod_5077_inner, "mod_5077");
    Operation_IFC mod_5078_inner <- mkRepeatStatic(8);
    Operation_IFC mod_5078 <- mkDebugOperation(mod_5078_inner, "mod_5078");
    Operation_IFC mod_5079_inner <- mkFlatten(1);
    Operation_IFC mod_5079 <- mkDebugOperation(mod_5079_inner, "mod_5079");
    Operation_IFC mod_5080_inner <- mkFlatten(0);
    Operation_IFC mod_5080 <- mkDebugOperation(mod_5080_inner, "mod_5080");
    Operation_IFC mod_5081_inner <- mkRepeatStatic(16);
    Operation_IFC mod_5081 <- mkDebugOperation(mod_5081_inner, "mod_5081");
    Operation_IFC mod_5082_inner <- mkRepeatStatic(2);
    Operation_IFC mod_5082 <- mkDebugOperation(mod_5082_inner, "mod_5082");
    PMU_IFC mod_5083_bufferize <- mkPMU(2);
    Operation_IFC mod_5083_inner = mod_5083_bufferize.operation;
    Operation_IFC mod_5083 <- mkDebugOperation(mod_5083_inner, "mod_5083");
    rule rule_6520;
        ChannelMessage t;
        t <- mod_5075.get(1);
        mod_5070.put(0, t);
    endrule
    rule rule_6521;
        ChannelMessage t;
        t <- mod_5058.get(0);
        mod_5062.put(0, t);
    endrule
    rule rule_6522;
        ChannelMessage t;
        t <- mod_5065.get(0);
        mod_5063.put(0, t);
    endrule
    rule rule_6523;
        ChannelMessage t;
        t <- mod_5074.get(0);
        mod_5073.put(0, t);
    endrule
    rule rule_6524;
        ChannelMessage t;
        t <- mod_5059.get(0);
        mod_5061.put(0, t);
    endrule
    rule rule_6525;
        ChannelMessage t;
        t <- mod_5047.get(0);
        mod_5083.put(0, t);
    endrule
    rule rule_6526;
        ChannelMessage t;
        t <- mod_5071.get(1);
        mod_5070.put(1, t);
    endrule
    rule rule_6527;
        ChannelMessage t;
        t <- mod_5072.get(0);
        mod_5071.put(1, t);
    endrule
    rule rule_6528;
        ChannelMessage t;
        t <- mod_5051.get(1);
        mod_5052.put(0, t);
    endrule
    rule rule_6529;
        ChannelMessage t;
        t <- mod_5082.get(0);
        mod_5049.put(1, t);
    endrule
    rule rule_6530;
        ChannelMessage t;
        t <- mod_5057.get(0);
        mod_5058.put(0, t);
    endrule
    rule rule_6531;
        ChannelMessage t;
        t <- mod_5073.get(0);
        mod_5071.put(0, t);
    endrule
    rule rule_6532;
        ChannelMessage t;
        t <- mod_5049.get(1);
        mod_5050.put(0, t);
    endrule
    rule rule_6533;
        ChannelMessage t;
        t <- mod_5055.get(0);
        mod_5067.put(0, t);
    endrule
    rule rule_6534;
        ChannelMessage t;
        t <- mod_5062.get(1);
        mod_5058.put(1, t);
    endrule
    rule rule_6535;
        ChannelMessage t;
        t <- mod_5083.get(0);
        mod_5083.put(1, t);
    endrule
    rule rule_6536;
        ChannelMessage t;
        t <- mod_5063.get(0);
        mod_5064.put(0, t);
    endrule
    rule rule_6537;
        ChannelMessage t;
        t <- mod_5050.get(1);
        mod_5051.put(0, t);
    endrule
    rule rule_6538;
        ChannelMessage t;
        t <- mod_5062.get(0);
        mod_5062.put(1, t);
    endrule
    rule rule_6539;
        ChannelMessage t;
        t <- mod_5080.get(0);
        mod_5079.put(0, t);
    endrule
    rule rule_6540;
        ChannelMessage t;
        t <- mod_5064.get(0);
        mod_5063.put(1, t);
    endrule
    rule rule_6541;
        ChannelMessage t;
        t <- mod_5067.get(0);
        mod_5055.put(1, t);
    endrule
    rule rule_6542;
        ChannelMessage t;
        t <- mod_5048.get(3);
        mod_5049.put(0, t);
    endrule
    rule rule_6543;
        ChannelMessage t;
        t <- mod_5077.get(1);
        mod_5052.put(1, t);
    endrule
    rule rule_6544;
        ChannelMessage t;
        t <- mod_5079.get(0);
        mod_5077.put(0, t);
    endrule
    rule rule_6545;
        ChannelMessage t;
        t <- mod_5071.get(0);
        mod_5072.put(0, t);
    endrule
    rule rule_6546;
        ChannelMessage t;
        t <- mod_5044.get(0);
        mod_5045.put(0, t);
    endrule
    rule rule_6547;
        ChannelMessage t;
        t <- mod_5045.get(0);
        mod_5046.put(0, t);
    endrule
    rule rule_6548;
        ChannelMessage t;
        t <- mod_5054.get(0);
        mod_5055.put(0, t);
    endrule
    rule rule_6549;
        ChannelMessage t;
        t <- mod_5055.get(1);
        mod_5056.put(0, t);
    endrule
    rule rule_6550;
        ChannelMessage t;
        t <- mod_5081.get(0);
        mod_5051.put(1, t);
    endrule
    rule rule_6551;
        ChannelMessage t;
        t <- mod_5061.get(1);
        mod_5059.put(1, t);
    endrule
    rule rule_6552;
        ChannelMessage t;
        t <- mod_5056.get(0);
        mod_5057.put(0, t);
    endrule
    rule rule_6553;
        ChannelMessage t;
        t <- mod_5058.get(1);
        mod_5059.put(0, t);
    endrule
    rule rule_6554;
        ChannelMessage t;
        t <- mod_5046.get(0);
        mod_5047.put(0, t);
    endrule
    rule rule_6555;
        ChannelMessage t;
        t <- mod_5070.get(0);
        mod_5069.put(0, t);
    endrule
    rule rule_6556;
        ChannelMessage t;
        t <- mod_5047.get(1);
        mod_5048.put(0, t);
    endrule
    rule rule_6557;
        ChannelMessage t;
        t <- mod_5059.get(1);
        mod_5060.put(1, t);
    endrule
    rule rule_6558;
        ChannelMessage t;
        t <- mod_5076.get(0);
        mod_5075.put(1, t);
    endrule
    rule rule_6559;
        ChannelMessage t;
        t <- mod_5078.get(0);
        mod_5077.put(1, t);
    endrule
    rule rule_6560;
        ChannelMessage t;
        t <- mod_5053.get(0);
        mod_5054.put(0, t);
    endrule
    rule rule_6561;
        ChannelMessage t;
        t <- mod_5077.get(0);
        mod_5078.put(0, t);
    endrule
    rule rule_6562;
        ChannelMessage t;
        t <- mod_5050.get(0);
        mod_5075.put(0, t);
    endrule
    rule rule_6563;
        ChannelMessage t;
        t <- mod_5052.get(0);
        mod_5053.put(0, t);
    endrule
    rule rule_6564;
        ChannelMessage t;
        t <- mod_5063.get(1);
        mod_5056.put(1, t);
    endrule
    rule rule_6565;
        ChannelMessage t;
        t <- mod_5051.get(0);
        mod_5081.put(0, t);
    endrule
    rule rule_6566;
        ChannelMessage t;
        t <- mod_5069.get(0);
        mod_5068.put(0, t);
    endrule
    rule rule_6567;
        ChannelMessage t;
        t <- mod_5083.get(1);
        mod_5047.put(1, t);
    endrule
    rule rule_6568;
        ChannelMessage t;
        t <- mod_5049.get(0);
        mod_5082.put(0, t);
    endrule
    rule rule_6569;
        ChannelMessage t;
        t <- mod_5061.get(0);
        mod_5061.put(1, t);
    endrule
    rule rule_6570;
        ChannelMessage t;
        t <- mod_5068.get(0);
        mod_5054.put(1, t);
    endrule
    rule rule_6571;
        ChannelMessage t;
        t <- mod_5066.get(0);
        mod_5065.put(0, t);
    endrule
    rule rule_6572;
        ChannelMessage t;
        t <- mod_5075.get(0);
        mod_5076.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_5044.put(0, t);
        end
        if (i == 1) begin
            mod_5060.put(0, t);
        end
        if (i == 2) begin
            mod_5066.put(0, t);
        end
        if (i == 3) begin
            mod_5074.put(0, t);
        end
        if (i == 4) begin
            mod_5080.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_5048.get(0);
        end
        if (i == 2) begin
            t <- mod_5048.get(1);
        end
        if (i == 3) begin
            t <- mod_5048.get(2);
        end
        if (i == 0) begin
            t <- mod_5060.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6158 (Operation_IFC);
    Operation_IFC mod_5085_inner <- mkReshape(2, 64);
    Operation_IFC mod_5085 <- mkDebugOperation(mod_5085_inner, "mod_5085");
    Operation_IFC mod_5086_inner <- mkFlatten(1);
    Operation_IFC mod_5086 <- mkDebugOperation(mod_5086_inner, "mod_5086");
    Operation_IFC mod_5087_inner <- mkFlatten(2);
    Operation_IFC mod_5087 <- mkDebugOperation(mod_5087_inner, "mod_5087");
    Operation_IFC mod_5088_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_5088 <- mkDebugOperation(mod_5088_inner, "mod_5088");
    Broadcast_IFC#(4) mod_5089_inner <- mkBroadcast(4);
    Operation_IFC mod_5089 <- mkDebugOperation(mod_5089_inner.op, "mod_5089");
    PMU_IFC mod_5090_bufferize <- mkPMU(2);
    Operation_IFC mod_5090_inner = mod_5090_bufferize.operation;
    Operation_IFC mod_5090 <- mkDebugOperation(mod_5090_inner, "mod_5090");
    Broadcast_IFC#(2) mod_5091_inner <- mkBroadcast(2);
    Operation_IFC mod_5091 <- mkDebugOperation(mod_5091_inner.op, "mod_5091");
    PMU_IFC mod_5092_bufferize <- mkPMU(1);
    Operation_IFC mod_5092_inner = mod_5092_bufferize.operation;
    Operation_IFC mod_5092 <- mkDebugOperation(mod_5092_inner, "mod_5092");
    Operation_IFC mod_5093_inner <- mkBinaryMap(1032, matmul_t_tile);
    Operation_IFC mod_5093 <- mkDebugOperation(mod_5093_inner, "mod_5093");
    Operation_IFC mod_5094_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_5094 <- mkDebugOperation(mod_5094_inner, "mod_5094");
    Operation_IFC mod_5095_inner <- mkBinaryMap(1800, mul_tile);
    Operation_IFC mod_5095 <- mkDebugOperation(mod_5095_inner, "mod_5095");
    PMU_IFC mod_5096_bufferize <- mkPMU(1);
    Operation_IFC mod_5096_inner = mod_5096_bufferize.operation;
    Operation_IFC mod_5096 <- mkDebugOperation(mod_5096_inner, "mod_5096");
    Operation_IFC mod_5097_inner <- mkBinaryMap(2315, matmul_t_tile);
    Operation_IFC mod_5097 <- mkDebugOperation(mod_5097_inner, "mod_5097");
    Operation_IFC mod_5098_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_5098 <- mkDebugOperation(mod_5098_inner, "mod_5098");
    Operation_IFC mod_5099_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_5099 <- mkDebugOperation(mod_5099_inner, "mod_5099");
    Operation_IFC mod_5100_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_5100 <- mkDebugOperation(mod_5100_inner, "mod_5100");
    Operation_IFC mod_5101_inner <- mkBinaryMap(2699, mul_tile);
    Operation_IFC mod_5101 <- mkDebugOperation(mod_5101_inner, "mod_5101");
    PMU_IFC mod_5102_bufferize <- mkPMU(1);
    Operation_IFC mod_5102_inner = mod_5102_bufferize.operation;
    Operation_IFC mod_5102 <- mkDebugOperation(mod_5102_inner, "mod_5102");
    PMU_IFC mod_5103_bufferize <- mkPMU(2);
    Operation_IFC mod_5103_inner = mod_5103_bufferize.operation;
    Operation_IFC mod_5103 <- mkDebugOperation(mod_5103_inner, "mod_5103");
    PMU_IFC mod_5104_bufferize <- mkPMU(2);
    Operation_IFC mod_5104_inner = mod_5104_bufferize.operation;
    Operation_IFC mod_5104 <- mkDebugOperation(mod_5104_inner, "mod_5104");
    Operation_IFC mod_5105_inner <- mkRepeatStatic(8);
    Operation_IFC mod_5105 <- mkDebugOperation(mod_5105_inner, "mod_5105");
    Operation_IFC mod_5106_inner <- mkFlatten(1);
    Operation_IFC mod_5106 <- mkDebugOperation(mod_5106_inner, "mod_5106");
    Operation_IFC mod_5107_inner <- mkFlatten(0);
    Operation_IFC mod_5107 <- mkDebugOperation(mod_5107_inner, "mod_5107");
    Operation_IFC mod_5108_inner <- mkRepeatStatic(3);
    Operation_IFC mod_5108 <- mkDebugOperation(mod_5108_inner, "mod_5108");
    Operation_IFC mod_5109_inner <- mkUnaryMap(1672, silu_tile);
    Operation_IFC mod_5109 <- mkDebugOperation(mod_5109_inner, "mod_5109");
    Operation_IFC mod_5110_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_5110 <- mkDebugOperation(mod_5110_inner, "mod_5110");
    Operation_IFC mod_5111_inner <- mkBinaryMap(1544, matmul_t_tile);
    Operation_IFC mod_5111 <- mkDebugOperation(mod_5111_inner, "mod_5111");
    PMU_IFC mod_5112_bufferize <- mkPMU(2);
    Operation_IFC mod_5112_inner = mod_5112_bufferize.operation;
    Operation_IFC mod_5112 <- mkDebugOperation(mod_5112_inner, "mod_5112");
    Operation_IFC mod_5113_inner <- mkRepeatStatic(8);
    Operation_IFC mod_5113 <- mkDebugOperation(mod_5113_inner, "mod_5113");
    Operation_IFC mod_5114_inner <- mkFlatten(1);
    Operation_IFC mod_5114 <- mkDebugOperation(mod_5114_inner, "mod_5114");
    Operation_IFC mod_5115_inner <- mkFlatten(0);
    Operation_IFC mod_5115 <- mkDebugOperation(mod_5115_inner, "mod_5115");
    PMU_IFC mod_5116_bufferize <- mkPMU(1);
    Operation_IFC mod_5116_inner = mod_5116_bufferize.operation;
    Operation_IFC mod_5116 <- mkDebugOperation(mod_5116_inner, "mod_5116");
    Operation_IFC mod_5117_inner <- mkRepeatStatic(16);
    Operation_IFC mod_5117 <- mkDebugOperation(mod_5117_inner, "mod_5117");
    PMU_IFC mod_5118_bufferize <- mkPMU(2);
    Operation_IFC mod_5118_inner = mod_5118_bufferize.operation;
    Operation_IFC mod_5118 <- mkDebugOperation(mod_5118_inner, "mod_5118");
    Operation_IFC mod_5119_inner <- mkRepeatStatic(8);
    Operation_IFC mod_5119 <- mkDebugOperation(mod_5119_inner, "mod_5119");
    Operation_IFC mod_5120_inner <- mkFlatten(1);
    Operation_IFC mod_5120 <- mkDebugOperation(mod_5120_inner, "mod_5120");
    Operation_IFC mod_5121_inner <- mkFlatten(0);
    Operation_IFC mod_5121 <- mkDebugOperation(mod_5121_inner, "mod_5121");
    Operation_IFC mod_5122_inner <- mkRepeatStatic(16);
    Operation_IFC mod_5122 <- mkDebugOperation(mod_5122_inner, "mod_5122");
    Operation_IFC mod_5123_inner <- mkRepeatStatic(2);
    Operation_IFC mod_5123 <- mkDebugOperation(mod_5123_inner, "mod_5123");
    PMU_IFC mod_5124_bufferize <- mkPMU(2);
    Operation_IFC mod_5124_inner = mod_5124_bufferize.operation;
    Operation_IFC mod_5124 <- mkDebugOperation(mod_5124_inner, "mod_5124");
    rule rule_6573;
        ChannelMessage t;
        t <- mod_5092.get(0);
        mod_5122.put(0, t);
    endrule
    rule rule_6574;
        ChannelMessage t;
        t <- mod_5090.get(1);
        mod_5091.put(0, t);
    endrule
    rule rule_6575;
        ChannelMessage t;
        t <- mod_5099.get(0);
        mod_5103.put(0, t);
    endrule
    rule rule_6576;
        ChannelMessage t;
        t <- mod_5116.get(0);
        mod_5117.put(0, t);
    endrule
    rule rule_6577;
        ChannelMessage t;
        t <- mod_5095.get(0);
        mod_5096.put(0, t);
    endrule
    rule rule_6578;
        ChannelMessage t;
        t <- mod_5115.get(0);
        mod_5114.put(0, t);
    endrule
    rule rule_6579;
        ChannelMessage t;
        t <- mod_5103.get(1);
        mod_5099.put(1, t);
    endrule
    rule rule_6580;
        ChannelMessage t;
        t <- mod_5088.get(0);
        mod_5124.put(0, t);
    endrule
    rule rule_6581;
        ChannelMessage t;
        t <- mod_5091.get(0);
        mod_5116.put(0, t);
    endrule
    rule rule_6582;
        ChannelMessage t;
        t <- mod_5104.get(1);
        mod_5097.put(1, t);
    endrule
    rule rule_6583;
        ChannelMessage t;
        t <- mod_5112.get(1);
        mod_5111.put(1, t);
    endrule
    rule rule_6584;
        ChannelMessage t;
        t <- mod_5099.get(1);
        mod_5100.put(0, t);
    endrule
    rule rule_6585;
        ChannelMessage t;
        t <- mod_5086.get(0);
        mod_5087.put(0, t);
    endrule
    rule rule_6586;
        ChannelMessage t;
        t <- mod_5122.get(0);
        mod_5092.put(1, t);
    endrule
    rule rule_6587;
        ChannelMessage t;
        t <- mod_5118.get(1);
        mod_5093.put(1, t);
    endrule
    rule rule_6588;
        ChannelMessage t;
        t <- mod_5113.get(0);
        mod_5112.put(1, t);
    endrule
    rule rule_6589;
        ChannelMessage t;
        t <- mod_5102.get(1);
        mod_5100.put(1, t);
    endrule
    rule rule_6590;
        ChannelMessage t;
        t <- mod_5109.get(0);
        mod_5095.put(1, t);
    endrule
    rule rule_6591;
        ChannelMessage t;
        t <- mod_5123.get(0);
        mod_5090.put(1, t);
    endrule
    rule rule_6592;
        ChannelMessage t;
        t <- mod_5090.get(0);
        mod_5123.put(0, t);
    endrule
    rule rule_6593;
        ChannelMessage t;
        t <- mod_5096.get(1);
        mod_5097.put(0, t);
    endrule
    rule rule_6594;
        ChannelMessage t;
        t <- mod_5108.get(0);
        mod_5096.put(1, t);
    endrule
    rule rule_6595;
        ChannelMessage t;
        t <- mod_5092.get(1);
        mod_5093.put(0, t);
    endrule
    rule rule_6596;
        ChannelMessage t;
        t <- mod_5085.get(0);
        mod_5086.put(0, t);
    endrule
    rule rule_6597;
        ChannelMessage t;
        t <- mod_5114.get(0);
        mod_5112.put(0, t);
    endrule
    rule rule_6598;
        ChannelMessage t;
        t <- mod_5116.get(1);
        mod_5111.put(0, t);
    endrule
    rule rule_6599;
        ChannelMessage t;
        t <- mod_5124.get(0);
        mod_5124.put(1, t);
    endrule
    rule rule_6600;
        ChannelMessage t;
        t <- mod_5100.get(0);
        mod_5102.put(0, t);
    endrule
    rule rule_6601;
        ChannelMessage t;
        t <- mod_5111.get(0);
        mod_5110.put(0, t);
    endrule
    rule rule_6602;
        ChannelMessage t;
        t <- mod_5100.get(1);
        mod_5101.put(1, t);
    endrule
    rule rule_6603;
        ChannelMessage t;
        t <- mod_5121.get(0);
        mod_5120.put(0, t);
    endrule
    rule rule_6604;
        ChannelMessage t;
        t <- mod_5087.get(0);
        mod_5088.put(0, t);
    endrule
    rule rule_6605;
        ChannelMessage t;
        t <- mod_5098.get(0);
        mod_5099.put(0, t);
    endrule
    rule rule_6606;
        ChannelMessage t;
        t <- mod_5118.get(0);
        mod_5119.put(0, t);
    endrule
    rule rule_6607;
        ChannelMessage t;
        t <- mod_5093.get(0);
        mod_5094.put(0, t);
    endrule
    rule rule_6608;
        ChannelMessage t;
        t <- mod_5104.get(0);
        mod_5105.put(0, t);
    endrule
    rule rule_6609;
        ChannelMessage t;
        t <- mod_5089.get(3);
        mod_5090.put(0, t);
    endrule
    rule rule_6610;
        ChannelMessage t;
        t <- mod_5096.get(0);
        mod_5108.put(0, t);
    endrule
    rule rule_6611;
        ChannelMessage t;
        t <- mod_5091.get(1);
        mod_5092.put(0, t);
    endrule
    rule rule_6612;
        ChannelMessage t;
        t <- mod_5107.get(0);
        mod_5106.put(0, t);
    endrule
    rule rule_6613;
        ChannelMessage t;
        t <- mod_5119.get(0);
        mod_5118.put(1, t);
    endrule
    rule rule_6614;
        ChannelMessage t;
        t <- mod_5110.get(0);
        mod_5109.put(0, t);
    endrule
    rule rule_6615;
        ChannelMessage t;
        t <- mod_5117.get(0);
        mod_5116.put(1, t);
    endrule
    rule rule_6616;
        ChannelMessage t;
        t <- mod_5112.get(0);
        mod_5113.put(0, t);
    endrule
    rule rule_6617;
        ChannelMessage t;
        t <- mod_5120.get(0);
        mod_5118.put(0, t);
    endrule
    rule rule_6618;
        ChannelMessage t;
        t <- mod_5097.get(0);
        mod_5098.put(0, t);
    endrule
    rule rule_6619;
        ChannelMessage t;
        t <- mod_5088.get(1);
        mod_5089.put(0, t);
    endrule
    rule rule_6620;
        ChannelMessage t;
        t <- mod_5103.get(0);
        mod_5103.put(1, t);
    endrule
    rule rule_6621;
        ChannelMessage t;
        t <- mod_5105.get(0);
        mod_5104.put(1, t);
    endrule
    rule rule_6622;
        ChannelMessage t;
        t <- mod_5124.get(1);
        mod_5088.put(1, t);
    endrule
    rule rule_6623;
        ChannelMessage t;
        t <- mod_5102.get(0);
        mod_5102.put(1, t);
    endrule
    rule rule_6624;
        ChannelMessage t;
        t <- mod_5106.get(0);
        mod_5104.put(0, t);
    endrule
    rule rule_6625;
        ChannelMessage t;
        t <- mod_5094.get(0);
        mod_5095.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_5085.put(0, t);
        end
        if (i == 1) begin
            mod_5101.put(0, t);
        end
        if (i == 2) begin
            mod_5107.put(0, t);
        end
        if (i == 3) begin
            mod_5115.put(0, t);
        end
        if (i == 4) begin
            mod_5121.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_5089.get(0);
        end
        if (i == 0) begin
            t <- mod_5089.get(1);
        end
        if (i == 1) begin
            t <- mod_5089.get(2);
        end
        if (i == 2) begin
            t <- mod_5101.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6159 (Operation_IFC);
    Operation_IFC mod_5126_inner <- mkReshape(2, 64);
    Operation_IFC mod_5126 <- mkDebugOperation(mod_5126_inner, "mod_5126");
    Operation_IFC mod_5127_inner <- mkFlatten(1);
    Operation_IFC mod_5127 <- mkDebugOperation(mod_5127_inner, "mod_5127");
    Operation_IFC mod_5128_inner <- mkFlatten(2);
    Operation_IFC mod_5128 <- mkDebugOperation(mod_5128_inner, "mod_5128");
    Operation_IFC mod_5129_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_5129 <- mkDebugOperation(mod_5129_inner, "mod_5129");
    Broadcast_IFC#(4) mod_5130_inner <- mkBroadcast(4);
    Operation_IFC mod_5130 <- mkDebugOperation(mod_5130_inner.op, "mod_5130");
    PMU_IFC mod_5131_bufferize <- mkPMU(2);
    Operation_IFC mod_5131_inner = mod_5131_bufferize.operation;
    Operation_IFC mod_5131 <- mkDebugOperation(mod_5131_inner, "mod_5131");
    Broadcast_IFC#(2) mod_5132_inner <- mkBroadcast(2);
    Operation_IFC mod_5132 <- mkDebugOperation(mod_5132_inner.op, "mod_5132");
    PMU_IFC mod_5133_bufferize <- mkPMU(1);
    Operation_IFC mod_5133_inner = mod_5133_bufferize.operation;
    Operation_IFC mod_5133 <- mkDebugOperation(mod_5133_inner, "mod_5133");
    Operation_IFC mod_5134_inner <- mkBinaryMap(1031, matmul_t_tile);
    Operation_IFC mod_5134 <- mkDebugOperation(mod_5134_inner, "mod_5134");
    Operation_IFC mod_5135_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_5135 <- mkDebugOperation(mod_5135_inner, "mod_5135");
    Operation_IFC mod_5136_inner <- mkBinaryMap(1799, mul_tile);
    Operation_IFC mod_5136 <- mkDebugOperation(mod_5136_inner, "mod_5136");
    PMU_IFC mod_5137_bufferize <- mkPMU(1);
    Operation_IFC mod_5137_inner = mod_5137_bufferize.operation;
    Operation_IFC mod_5137 <- mkDebugOperation(mod_5137_inner, "mod_5137");
    Operation_IFC mod_5138_inner <- mkBinaryMap(2313, matmul_t_tile);
    Operation_IFC mod_5138 <- mkDebugOperation(mod_5138_inner, "mod_5138");
    Operation_IFC mod_5139_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_5139 <- mkDebugOperation(mod_5139_inner, "mod_5139");
    Operation_IFC mod_5140_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_5140 <- mkDebugOperation(mod_5140_inner, "mod_5140");
    Operation_IFC mod_5141_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_5141 <- mkDebugOperation(mod_5141_inner, "mod_5141");
    Operation_IFC mod_5142_inner <- mkBinaryMap(2698, mul_tile);
    Operation_IFC mod_5142 <- mkDebugOperation(mod_5142_inner, "mod_5142");
    PMU_IFC mod_5143_bufferize <- mkPMU(1);
    Operation_IFC mod_5143_inner = mod_5143_bufferize.operation;
    Operation_IFC mod_5143 <- mkDebugOperation(mod_5143_inner, "mod_5143");
    PMU_IFC mod_5144_bufferize <- mkPMU(2);
    Operation_IFC mod_5144_inner = mod_5144_bufferize.operation;
    Operation_IFC mod_5144 <- mkDebugOperation(mod_5144_inner, "mod_5144");
    PMU_IFC mod_5145_bufferize <- mkPMU(2);
    Operation_IFC mod_5145_inner = mod_5145_bufferize.operation;
    Operation_IFC mod_5145 <- mkDebugOperation(mod_5145_inner, "mod_5145");
    Operation_IFC mod_5146_inner <- mkRepeatStatic(8);
    Operation_IFC mod_5146 <- mkDebugOperation(mod_5146_inner, "mod_5146");
    Operation_IFC mod_5147_inner <- mkFlatten(1);
    Operation_IFC mod_5147 <- mkDebugOperation(mod_5147_inner, "mod_5147");
    Operation_IFC mod_5148_inner <- mkFlatten(0);
    Operation_IFC mod_5148 <- mkDebugOperation(mod_5148_inner, "mod_5148");
    Operation_IFC mod_5149_inner <- mkRepeatStatic(3);
    Operation_IFC mod_5149 <- mkDebugOperation(mod_5149_inner, "mod_5149");
    Operation_IFC mod_5150_inner <- mkUnaryMap(1671, silu_tile);
    Operation_IFC mod_5150 <- mkDebugOperation(mod_5150_inner, "mod_5150");
    Operation_IFC mod_5151_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_5151 <- mkDebugOperation(mod_5151_inner, "mod_5151");
    Operation_IFC mod_5152_inner <- mkBinaryMap(1543, matmul_t_tile);
    Operation_IFC mod_5152 <- mkDebugOperation(mod_5152_inner, "mod_5152");
    PMU_IFC mod_5153_bufferize <- mkPMU(2);
    Operation_IFC mod_5153_inner = mod_5153_bufferize.operation;
    Operation_IFC mod_5153 <- mkDebugOperation(mod_5153_inner, "mod_5153");
    Operation_IFC mod_5154_inner <- mkRepeatStatic(8);
    Operation_IFC mod_5154 <- mkDebugOperation(mod_5154_inner, "mod_5154");
    Operation_IFC mod_5155_inner <- mkFlatten(1);
    Operation_IFC mod_5155 <- mkDebugOperation(mod_5155_inner, "mod_5155");
    Operation_IFC mod_5156_inner <- mkFlatten(0);
    Operation_IFC mod_5156 <- mkDebugOperation(mod_5156_inner, "mod_5156");
    PMU_IFC mod_5157_bufferize <- mkPMU(1);
    Operation_IFC mod_5157_inner = mod_5157_bufferize.operation;
    Operation_IFC mod_5157 <- mkDebugOperation(mod_5157_inner, "mod_5157");
    Operation_IFC mod_5158_inner <- mkRepeatStatic(16);
    Operation_IFC mod_5158 <- mkDebugOperation(mod_5158_inner, "mod_5158");
    PMU_IFC mod_5159_bufferize <- mkPMU(2);
    Operation_IFC mod_5159_inner = mod_5159_bufferize.operation;
    Operation_IFC mod_5159 <- mkDebugOperation(mod_5159_inner, "mod_5159");
    Operation_IFC mod_5160_inner <- mkRepeatStatic(8);
    Operation_IFC mod_5160 <- mkDebugOperation(mod_5160_inner, "mod_5160");
    Operation_IFC mod_5161_inner <- mkFlatten(1);
    Operation_IFC mod_5161 <- mkDebugOperation(mod_5161_inner, "mod_5161");
    Operation_IFC mod_5162_inner <- mkFlatten(0);
    Operation_IFC mod_5162 <- mkDebugOperation(mod_5162_inner, "mod_5162");
    Operation_IFC mod_5163_inner <- mkRepeatStatic(16);
    Operation_IFC mod_5163 <- mkDebugOperation(mod_5163_inner, "mod_5163");
    Operation_IFC mod_5164_inner <- mkRepeatStatic(2);
    Operation_IFC mod_5164 <- mkDebugOperation(mod_5164_inner, "mod_5164");
    PMU_IFC mod_5165_bufferize <- mkPMU(2);
    Operation_IFC mod_5165_inner = mod_5165_bufferize.operation;
    Operation_IFC mod_5165 <- mkDebugOperation(mod_5165_inner, "mod_5165");
    rule rule_6626;
        ChannelMessage t;
        t <- mod_5138.get(0);
        mod_5139.put(0, t);
    endrule
    rule rule_6627;
        ChannelMessage t;
        t <- mod_5154.get(0);
        mod_5153.put(1, t);
    endrule
    rule rule_6628;
        ChannelMessage t;
        t <- mod_5150.get(0);
        mod_5136.put(1, t);
    endrule
    rule rule_6629;
        ChannelMessage t;
        t <- mod_5160.get(0);
        mod_5159.put(1, t);
    endrule
    rule rule_6630;
        ChannelMessage t;
        t <- mod_5129.get(0);
        mod_5165.put(0, t);
    endrule
    rule rule_6631;
        ChannelMessage t;
        t <- mod_5153.get(0);
        mod_5154.put(0, t);
    endrule
    rule rule_6632;
        ChannelMessage t;
        t <- mod_5157.get(0);
        mod_5158.put(0, t);
    endrule
    rule rule_6633;
        ChannelMessage t;
        t <- mod_5158.get(0);
        mod_5157.put(1, t);
    endrule
    rule rule_6634;
        ChannelMessage t;
        t <- mod_5159.get(1);
        mod_5134.put(1, t);
    endrule
    rule rule_6635;
        ChannelMessage t;
        t <- mod_5140.get(1);
        mod_5141.put(0, t);
    endrule
    rule rule_6636;
        ChannelMessage t;
        t <- mod_5131.get(0);
        mod_5164.put(0, t);
    endrule
    rule rule_6637;
        ChannelMessage t;
        t <- mod_5140.get(0);
        mod_5144.put(0, t);
    endrule
    rule rule_6638;
        ChannelMessage t;
        t <- mod_5151.get(0);
        mod_5150.put(0, t);
    endrule
    rule rule_6639;
        ChannelMessage t;
        t <- mod_5126.get(0);
        mod_5127.put(0, t);
    endrule
    rule rule_6640;
        ChannelMessage t;
        t <- mod_5152.get(0);
        mod_5151.put(0, t);
    endrule
    rule rule_6641;
        ChannelMessage t;
        t <- mod_5149.get(0);
        mod_5137.put(1, t);
    endrule
    rule rule_6642;
        ChannelMessage t;
        t <- mod_5133.get(1);
        mod_5134.put(0, t);
    endrule
    rule rule_6643;
        ChannelMessage t;
        t <- mod_5132.get(1);
        mod_5133.put(0, t);
    endrule
    rule rule_6644;
        ChannelMessage t;
        t <- mod_5153.get(1);
        mod_5152.put(1, t);
    endrule
    rule rule_6645;
        ChannelMessage t;
        t <- mod_5143.get(1);
        mod_5141.put(1, t);
    endrule
    rule rule_6646;
        ChannelMessage t;
        t <- mod_5147.get(0);
        mod_5145.put(0, t);
    endrule
    rule rule_6647;
        ChannelMessage t;
        t <- mod_5139.get(0);
        mod_5140.put(0, t);
    endrule
    rule rule_6648;
        ChannelMessage t;
        t <- mod_5144.get(0);
        mod_5144.put(1, t);
    endrule
    rule rule_6649;
        ChannelMessage t;
        t <- mod_5143.get(0);
        mod_5143.put(1, t);
    endrule
    rule rule_6650;
        ChannelMessage t;
        t <- mod_5148.get(0);
        mod_5147.put(0, t);
    endrule
    rule rule_6651;
        ChannelMessage t;
        t <- mod_5155.get(0);
        mod_5153.put(0, t);
    endrule
    rule rule_6652;
        ChannelMessage t;
        t <- mod_5128.get(0);
        mod_5129.put(0, t);
    endrule
    rule rule_6653;
        ChannelMessage t;
        t <- mod_5162.get(0);
        mod_5161.put(0, t);
    endrule
    rule rule_6654;
        ChannelMessage t;
        t <- mod_5144.get(1);
        mod_5140.put(1, t);
    endrule
    rule rule_6655;
        ChannelMessage t;
        t <- mod_5146.get(0);
        mod_5145.put(1, t);
    endrule
    rule rule_6656;
        ChannelMessage t;
        t <- mod_5145.get(0);
        mod_5146.put(0, t);
    endrule
    rule rule_6657;
        ChannelMessage t;
        t <- mod_5165.get(1);
        mod_5129.put(1, t);
    endrule
    rule rule_6658;
        ChannelMessage t;
        t <- mod_5137.get(0);
        mod_5149.put(0, t);
    endrule
    rule rule_6659;
        ChannelMessage t;
        t <- mod_5133.get(0);
        mod_5163.put(0, t);
    endrule
    rule rule_6660;
        ChannelMessage t;
        t <- mod_5134.get(0);
        mod_5135.put(0, t);
    endrule
    rule rule_6661;
        ChannelMessage t;
        t <- mod_5164.get(0);
        mod_5131.put(1, t);
    endrule
    rule rule_6662;
        ChannelMessage t;
        t <- mod_5129.get(1);
        mod_5130.put(0, t);
    endrule
    rule rule_6663;
        ChannelMessage t;
        t <- mod_5130.get(3);
        mod_5131.put(0, t);
    endrule
    rule rule_6664;
        ChannelMessage t;
        t <- mod_5136.get(0);
        mod_5137.put(0, t);
    endrule
    rule rule_6665;
        ChannelMessage t;
        t <- mod_5145.get(1);
        mod_5138.put(1, t);
    endrule
    rule rule_6666;
        ChannelMessage t;
        t <- mod_5157.get(1);
        mod_5152.put(0, t);
    endrule
    rule rule_6667;
        ChannelMessage t;
        t <- mod_5161.get(0);
        mod_5159.put(0, t);
    endrule
    rule rule_6668;
        ChannelMessage t;
        t <- mod_5165.get(0);
        mod_5165.put(1, t);
    endrule
    rule rule_6669;
        ChannelMessage t;
        t <- mod_5137.get(1);
        mod_5138.put(0, t);
    endrule
    rule rule_6670;
        ChannelMessage t;
        t <- mod_5156.get(0);
        mod_5155.put(0, t);
    endrule
    rule rule_6671;
        ChannelMessage t;
        t <- mod_5159.get(0);
        mod_5160.put(0, t);
    endrule
    rule rule_6672;
        ChannelMessage t;
        t <- mod_5132.get(0);
        mod_5157.put(0, t);
    endrule
    rule rule_6673;
        ChannelMessage t;
        t <- mod_5141.get(1);
        mod_5142.put(1, t);
    endrule
    rule rule_6674;
        ChannelMessage t;
        t <- mod_5127.get(0);
        mod_5128.put(0, t);
    endrule
    rule rule_6675;
        ChannelMessage t;
        t <- mod_5141.get(0);
        mod_5143.put(0, t);
    endrule
    rule rule_6676;
        ChannelMessage t;
        t <- mod_5163.get(0);
        mod_5133.put(1, t);
    endrule
    rule rule_6677;
        ChannelMessage t;
        t <- mod_5131.get(1);
        mod_5132.put(0, t);
    endrule
    rule rule_6678;
        ChannelMessage t;
        t <- mod_5135.get(0);
        mod_5136.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_5126.put(0, t);
        end
        if (i == 1) begin
            mod_5142.put(0, t);
        end
        if (i == 2) begin
            mod_5148.put(0, t);
        end
        if (i == 3) begin
            mod_5156.put(0, t);
        end
        if (i == 4) begin
            mod_5162.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 3) begin
            t <- mod_5130.get(0);
        end
        if (i == 0) begin
            t <- mod_5130.get(1);
        end
        if (i == 2) begin
            t <- mod_5130.get(2);
        end
        if (i == 1) begin
            t <- mod_5142.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6160 (Operation_IFC);
    Operation_IFC mod_5167_inner <- mkReshape(2, 64);
    Operation_IFC mod_5167 <- mkDebugOperation(mod_5167_inner, "mod_5167");
    Operation_IFC mod_5168_inner <- mkFlatten(1);
    Operation_IFC mod_5168 <- mkDebugOperation(mod_5168_inner, "mod_5168");
    Operation_IFC mod_5169_inner <- mkFlatten(2);
    Operation_IFC mod_5169 <- mkDebugOperation(mod_5169_inner, "mod_5169");
    Operation_IFC mod_5170_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_5170 <- mkDebugOperation(mod_5170_inner, "mod_5170");
    Broadcast_IFC#(4) mod_5171_inner <- mkBroadcast(4);
    Operation_IFC mod_5171 <- mkDebugOperation(mod_5171_inner.op, "mod_5171");
    PMU_IFC mod_5172_bufferize <- mkPMU(2);
    Operation_IFC mod_5172_inner = mod_5172_bufferize.operation;
    Operation_IFC mod_5172 <- mkDebugOperation(mod_5172_inner, "mod_5172");
    Broadcast_IFC#(2) mod_5173_inner <- mkBroadcast(2);
    Operation_IFC mod_5173 <- mkDebugOperation(mod_5173_inner.op, "mod_5173");
    PMU_IFC mod_5174_bufferize <- mkPMU(1);
    Operation_IFC mod_5174_inner = mod_5174_bufferize.operation;
    Operation_IFC mod_5174 <- mkDebugOperation(mod_5174_inner, "mod_5174");
    Operation_IFC mod_5175_inner <- mkBinaryMap(1030, matmul_t_tile);
    Operation_IFC mod_5175 <- mkDebugOperation(mod_5175_inner, "mod_5175");
    Operation_IFC mod_5176_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_5176 <- mkDebugOperation(mod_5176_inner, "mod_5176");
    Operation_IFC mod_5177_inner <- mkBinaryMap(1798, mul_tile);
    Operation_IFC mod_5177 <- mkDebugOperation(mod_5177_inner, "mod_5177");
    PMU_IFC mod_5178_bufferize <- mkPMU(1);
    Operation_IFC mod_5178_inner = mod_5178_bufferize.operation;
    Operation_IFC mod_5178 <- mkDebugOperation(mod_5178_inner, "mod_5178");
    Operation_IFC mod_5179_inner <- mkBinaryMap(2311, matmul_t_tile);
    Operation_IFC mod_5179 <- mkDebugOperation(mod_5179_inner, "mod_5179");
    Operation_IFC mod_5180_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_5180 <- mkDebugOperation(mod_5180_inner, "mod_5180");
    Operation_IFC mod_5181_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_5181 <- mkDebugOperation(mod_5181_inner, "mod_5181");
    Operation_IFC mod_5182_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_5182 <- mkDebugOperation(mod_5182_inner, "mod_5182");
    Operation_IFC mod_5183_inner <- mkBinaryMap(2697, mul_tile);
    Operation_IFC mod_5183 <- mkDebugOperation(mod_5183_inner, "mod_5183");
    PMU_IFC mod_5184_bufferize <- mkPMU(1);
    Operation_IFC mod_5184_inner = mod_5184_bufferize.operation;
    Operation_IFC mod_5184 <- mkDebugOperation(mod_5184_inner, "mod_5184");
    PMU_IFC mod_5185_bufferize <- mkPMU(2);
    Operation_IFC mod_5185_inner = mod_5185_bufferize.operation;
    Operation_IFC mod_5185 <- mkDebugOperation(mod_5185_inner, "mod_5185");
    PMU_IFC mod_5186_bufferize <- mkPMU(2);
    Operation_IFC mod_5186_inner = mod_5186_bufferize.operation;
    Operation_IFC mod_5186 <- mkDebugOperation(mod_5186_inner, "mod_5186");
    Operation_IFC mod_5187_inner <- mkRepeatStatic(8);
    Operation_IFC mod_5187 <- mkDebugOperation(mod_5187_inner, "mod_5187");
    Operation_IFC mod_5188_inner <- mkFlatten(1);
    Operation_IFC mod_5188 <- mkDebugOperation(mod_5188_inner, "mod_5188");
    Operation_IFC mod_5189_inner <- mkFlatten(0);
    Operation_IFC mod_5189 <- mkDebugOperation(mod_5189_inner, "mod_5189");
    Operation_IFC mod_5190_inner <- mkRepeatStatic(3);
    Operation_IFC mod_5190 <- mkDebugOperation(mod_5190_inner, "mod_5190");
    Operation_IFC mod_5191_inner <- mkUnaryMap(1670, silu_tile);
    Operation_IFC mod_5191 <- mkDebugOperation(mod_5191_inner, "mod_5191");
    Operation_IFC mod_5192_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_5192 <- mkDebugOperation(mod_5192_inner, "mod_5192");
    Operation_IFC mod_5193_inner <- mkBinaryMap(1542, matmul_t_tile);
    Operation_IFC mod_5193 <- mkDebugOperation(mod_5193_inner, "mod_5193");
    PMU_IFC mod_5194_bufferize <- mkPMU(2);
    Operation_IFC mod_5194_inner = mod_5194_bufferize.operation;
    Operation_IFC mod_5194 <- mkDebugOperation(mod_5194_inner, "mod_5194");
    Operation_IFC mod_5195_inner <- mkRepeatStatic(8);
    Operation_IFC mod_5195 <- mkDebugOperation(mod_5195_inner, "mod_5195");
    Operation_IFC mod_5196_inner <- mkFlatten(1);
    Operation_IFC mod_5196 <- mkDebugOperation(mod_5196_inner, "mod_5196");
    Operation_IFC mod_5197_inner <- mkFlatten(0);
    Operation_IFC mod_5197 <- mkDebugOperation(mod_5197_inner, "mod_5197");
    PMU_IFC mod_5198_bufferize <- mkPMU(1);
    Operation_IFC mod_5198_inner = mod_5198_bufferize.operation;
    Operation_IFC mod_5198 <- mkDebugOperation(mod_5198_inner, "mod_5198");
    Operation_IFC mod_5199_inner <- mkRepeatStatic(16);
    Operation_IFC mod_5199 <- mkDebugOperation(mod_5199_inner, "mod_5199");
    PMU_IFC mod_5200_bufferize <- mkPMU(2);
    Operation_IFC mod_5200_inner = mod_5200_bufferize.operation;
    Operation_IFC mod_5200 <- mkDebugOperation(mod_5200_inner, "mod_5200");
    Operation_IFC mod_5201_inner <- mkRepeatStatic(8);
    Operation_IFC mod_5201 <- mkDebugOperation(mod_5201_inner, "mod_5201");
    Operation_IFC mod_5202_inner <- mkFlatten(1);
    Operation_IFC mod_5202 <- mkDebugOperation(mod_5202_inner, "mod_5202");
    Operation_IFC mod_5203_inner <- mkFlatten(0);
    Operation_IFC mod_5203 <- mkDebugOperation(mod_5203_inner, "mod_5203");
    Operation_IFC mod_5204_inner <- mkRepeatStatic(16);
    Operation_IFC mod_5204 <- mkDebugOperation(mod_5204_inner, "mod_5204");
    Operation_IFC mod_5205_inner <- mkRepeatStatic(2);
    Operation_IFC mod_5205 <- mkDebugOperation(mod_5205_inner, "mod_5205");
    PMU_IFC mod_5206_bufferize <- mkPMU(2);
    Operation_IFC mod_5206_inner = mod_5206_bufferize.operation;
    Operation_IFC mod_5206 <- mkDebugOperation(mod_5206_inner, "mod_5206");
    rule rule_6679;
        ChannelMessage t;
        t <- mod_5174.get(0);
        mod_5204.put(0, t);
    endrule
    rule rule_6680;
        ChannelMessage t;
        t <- mod_5182.get(1);
        mod_5183.put(1, t);
    endrule
    rule rule_6681;
        ChannelMessage t;
        t <- mod_5197.get(0);
        mod_5196.put(0, t);
    endrule
    rule rule_6682;
        ChannelMessage t;
        t <- mod_5200.get(0);
        mod_5201.put(0, t);
    endrule
    rule rule_6683;
        ChannelMessage t;
        t <- mod_5168.get(0);
        mod_5169.put(0, t);
    endrule
    rule rule_6684;
        ChannelMessage t;
        t <- mod_5181.get(1);
        mod_5182.put(0, t);
    endrule
    rule rule_6685;
        ChannelMessage t;
        t <- mod_5184.get(0);
        mod_5184.put(1, t);
    endrule
    rule rule_6686;
        ChannelMessage t;
        t <- mod_5182.get(0);
        mod_5184.put(0, t);
    endrule
    rule rule_6687;
        ChannelMessage t;
        t <- mod_5173.get(1);
        mod_5174.put(0, t);
    endrule
    rule rule_6688;
        ChannelMessage t;
        t <- mod_5191.get(0);
        mod_5177.put(1, t);
    endrule
    rule rule_6689;
        ChannelMessage t;
        t <- mod_5167.get(0);
        mod_5168.put(0, t);
    endrule
    rule rule_6690;
        ChannelMessage t;
        t <- mod_5180.get(0);
        mod_5181.put(0, t);
    endrule
    rule rule_6691;
        ChannelMessage t;
        t <- mod_5186.get(0);
        mod_5187.put(0, t);
    endrule
    rule rule_6692;
        ChannelMessage t;
        t <- mod_5203.get(0);
        mod_5202.put(0, t);
    endrule
    rule rule_6693;
        ChannelMessage t;
        t <- mod_5170.get(0);
        mod_5206.put(0, t);
    endrule
    rule rule_6694;
        ChannelMessage t;
        t <- mod_5184.get(1);
        mod_5182.put(1, t);
    endrule
    rule rule_6695;
        ChannelMessage t;
        t <- mod_5190.get(0);
        mod_5178.put(1, t);
    endrule
    rule rule_6696;
        ChannelMessage t;
        t <- mod_5196.get(0);
        mod_5194.put(0, t);
    endrule
    rule rule_6697;
        ChannelMessage t;
        t <- mod_5198.get(0);
        mod_5199.put(0, t);
    endrule
    rule rule_6698;
        ChannelMessage t;
        t <- mod_5169.get(0);
        mod_5170.put(0, t);
    endrule
    rule rule_6699;
        ChannelMessage t;
        t <- mod_5179.get(0);
        mod_5180.put(0, t);
    endrule
    rule rule_6700;
        ChannelMessage t;
        t <- mod_5205.get(0);
        mod_5172.put(1, t);
    endrule
    rule rule_6701;
        ChannelMessage t;
        t <- mod_5170.get(1);
        mod_5171.put(0, t);
    endrule
    rule rule_6702;
        ChannelMessage t;
        t <- mod_5204.get(0);
        mod_5174.put(1, t);
    endrule
    rule rule_6703;
        ChannelMessage t;
        t <- mod_5193.get(0);
        mod_5192.put(0, t);
    endrule
    rule rule_6704;
        ChannelMessage t;
        t <- mod_5187.get(0);
        mod_5186.put(1, t);
    endrule
    rule rule_6705;
        ChannelMessage t;
        t <- mod_5185.get(1);
        mod_5181.put(1, t);
    endrule
    rule rule_6706;
        ChannelMessage t;
        t <- mod_5198.get(1);
        mod_5193.put(0, t);
    endrule
    rule rule_6707;
        ChannelMessage t;
        t <- mod_5202.get(0);
        mod_5200.put(0, t);
    endrule
    rule rule_6708;
        ChannelMessage t;
        t <- mod_5178.get(1);
        mod_5179.put(0, t);
    endrule
    rule rule_6709;
        ChannelMessage t;
        t <- mod_5171.get(3);
        mod_5172.put(0, t);
    endrule
    rule rule_6710;
        ChannelMessage t;
        t <- mod_5173.get(0);
        mod_5198.put(0, t);
    endrule
    rule rule_6711;
        ChannelMessage t;
        t <- mod_5185.get(0);
        mod_5185.put(1, t);
    endrule
    rule rule_6712;
        ChannelMessage t;
        t <- mod_5174.get(1);
        mod_5175.put(0, t);
    endrule
    rule rule_6713;
        ChannelMessage t;
        t <- mod_5172.get(1);
        mod_5173.put(0, t);
    endrule
    rule rule_6714;
        ChannelMessage t;
        t <- mod_5175.get(0);
        mod_5176.put(0, t);
    endrule
    rule rule_6715;
        ChannelMessage t;
        t <- mod_5192.get(0);
        mod_5191.put(0, t);
    endrule
    rule rule_6716;
        ChannelMessage t;
        t <- mod_5199.get(0);
        mod_5198.put(1, t);
    endrule
    rule rule_6717;
        ChannelMessage t;
        t <- mod_5206.get(1);
        mod_5170.put(1, t);
    endrule
    rule rule_6718;
        ChannelMessage t;
        t <- mod_5195.get(0);
        mod_5194.put(1, t);
    endrule
    rule rule_6719;
        ChannelMessage t;
        t <- mod_5177.get(0);
        mod_5178.put(0, t);
    endrule
    rule rule_6720;
        ChannelMessage t;
        t <- mod_5206.get(0);
        mod_5206.put(1, t);
    endrule
    rule rule_6721;
        ChannelMessage t;
        t <- mod_5181.get(0);
        mod_5185.put(0, t);
    endrule
    rule rule_6722;
        ChannelMessage t;
        t <- mod_5188.get(0);
        mod_5186.put(0, t);
    endrule
    rule rule_6723;
        ChannelMessage t;
        t <- mod_5186.get(1);
        mod_5179.put(1, t);
    endrule
    rule rule_6724;
        ChannelMessage t;
        t <- mod_5176.get(0);
        mod_5177.put(0, t);
    endrule
    rule rule_6725;
        ChannelMessage t;
        t <- mod_5178.get(0);
        mod_5190.put(0, t);
    endrule
    rule rule_6726;
        ChannelMessage t;
        t <- mod_5172.get(0);
        mod_5205.put(0, t);
    endrule
    rule rule_6727;
        ChannelMessage t;
        t <- mod_5200.get(1);
        mod_5175.put(1, t);
    endrule
    rule rule_6728;
        ChannelMessage t;
        t <- mod_5194.get(1);
        mod_5193.put(1, t);
    endrule
    rule rule_6729;
        ChannelMessage t;
        t <- mod_5189.get(0);
        mod_5188.put(0, t);
    endrule
    rule rule_6730;
        ChannelMessage t;
        t <- mod_5194.get(0);
        mod_5195.put(0, t);
    endrule
    rule rule_6731;
        ChannelMessage t;
        t <- mod_5201.get(0);
        mod_5200.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_5167.put(0, t);
        end
        if (i == 1) begin
            mod_5183.put(0, t);
        end
        if (i == 2) begin
            mod_5189.put(0, t);
        end
        if (i == 3) begin
            mod_5197.put(0, t);
        end
        if (i == 4) begin
            mod_5203.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_5171.get(0);
        end
        if (i == 3) begin
            t <- mod_5171.get(1);
        end
        if (i == 0) begin
            t <- mod_5171.get(2);
        end
        if (i == 2) begin
            t <- mod_5183.get(0);
        end

        return t;
    endmethod
endmodule
(* synthesize *)
module mkHypernode_6161 (Operation_IFC);
    Operation_IFC mod_5208_inner <- mkReshape(2, 64);
    Operation_IFC mod_5208 <- mkDebugOperation(mod_5208_inner, "mod_5208");
    Operation_IFC mod_5209_inner <- mkFlatten(1);
    Operation_IFC mod_5209 <- mkDebugOperation(mod_5209_inner, "mod_5209");
    Operation_IFC mod_5210_inner <- mkFlatten(2);
    Operation_IFC mod_5210 <- mkDebugOperation(mod_5210_inner, "mod_5210");
    Operation_IFC mod_5211_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_5211 <- mkDebugOperation(mod_5211_inner, "mod_5211");
    Broadcast_IFC#(4) mod_5212_inner <- mkBroadcast(4);
    Operation_IFC mod_5212 <- mkDebugOperation(mod_5212_inner.op, "mod_5212");
    PMU_IFC mod_5213_bufferize <- mkPMU(2);
    Operation_IFC mod_5213_inner = mod_5213_bufferize.operation;
    Operation_IFC mod_5213 <- mkDebugOperation(mod_5213_inner, "mod_5213");
    Broadcast_IFC#(2) mod_5214_inner <- mkBroadcast(2);
    Operation_IFC mod_5214 <- mkDebugOperation(mod_5214_inner.op, "mod_5214");
    PMU_IFC mod_5215_bufferize <- mkPMU(1);
    Operation_IFC mod_5215_inner = mod_5215_bufferize.operation;
    Operation_IFC mod_5215 <- mkDebugOperation(mod_5215_inner, "mod_5215");
    Operation_IFC mod_5216_inner <- mkBinaryMap(1029, matmul_t_tile);
    Operation_IFC mod_5216 <- mkDebugOperation(mod_5216_inner, "mod_5216");
    Operation_IFC mod_5217_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_5217 <- mkDebugOperation(mod_5217_inner, "mod_5217");
    Operation_IFC mod_5218_inner <- mkBinaryMap(1797, mul_tile);
    Operation_IFC mod_5218 <- mkDebugOperation(mod_5218_inner, "mod_5218");
    PMU_IFC mod_5219_bufferize <- mkPMU(1);
    Operation_IFC mod_5219_inner = mod_5219_bufferize.operation;
    Operation_IFC mod_5219 <- mkDebugOperation(mod_5219_inner, "mod_5219");
    Operation_IFC mod_5220_inner <- mkBinaryMap(2309, matmul_t_tile);
    Operation_IFC mod_5220 <- mkDebugOperation(mod_5220_inner, "mod_5220");
    Operation_IFC mod_5221_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_5221 <- mkDebugOperation(mod_5221_inner, "mod_5221");
    Operation_IFC mod_5222_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_5222 <- mkDebugOperation(mod_5222_inner, "mod_5222");
    Operation_IFC mod_5223_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_5223 <- mkDebugOperation(mod_5223_inner, "mod_5223");
    Operation_IFC mod_5224_inner <- mkBinaryMap(2696, mul_tile);
    Operation_IFC mod_5224 <- mkDebugOperation(mod_5224_inner, "mod_5224");
    PMU_IFC mod_5225_bufferize <- mkPMU(1);
    Operation_IFC mod_5225_inner = mod_5225_bufferize.operation;
    Operation_IFC mod_5225 <- mkDebugOperation(mod_5225_inner, "mod_5225");
    PMU_IFC mod_5226_bufferize <- mkPMU(2);
    Operation_IFC mod_5226_inner = mod_5226_bufferize.operation;
    Operation_IFC mod_5226 <- mkDebugOperation(mod_5226_inner, "mod_5226");
    PMU_IFC mod_5227_bufferize <- mkPMU(2);
    Operation_IFC mod_5227_inner = mod_5227_bufferize.operation;
    Operation_IFC mod_5227 <- mkDebugOperation(mod_5227_inner, "mod_5227");
    Operation_IFC mod_5228_inner <- mkRepeatStatic(8);
    Operation_IFC mod_5228 <- mkDebugOperation(mod_5228_inner, "mod_5228");
    Operation_IFC mod_5229_inner <- mkFlatten(1);
    Operation_IFC mod_5229 <- mkDebugOperation(mod_5229_inner, "mod_5229");
    Operation_IFC mod_5230_inner <- mkFlatten(0);
    Operation_IFC mod_5230 <- mkDebugOperation(mod_5230_inner, "mod_5230");
    Operation_IFC mod_5231_inner <- mkRepeatStatic(3);
    Operation_IFC mod_5231 <- mkDebugOperation(mod_5231_inner, "mod_5231");
    Operation_IFC mod_5232_inner <- mkUnaryMap(1669, silu_tile);
    Operation_IFC mod_5232 <- mkDebugOperation(mod_5232_inner, "mod_5232");
    Operation_IFC mod_5233_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_5233 <- mkDebugOperation(mod_5233_inner, "mod_5233");
    Operation_IFC mod_5234_inner <- mkBinaryMap(1541, matmul_t_tile);
    Operation_IFC mod_5234 <- mkDebugOperation(mod_5234_inner, "mod_5234");
    PMU_IFC mod_5235_bufferize <- mkPMU(2);
    Operation_IFC mod_5235_inner = mod_5235_bufferize.operation;
    Operation_IFC mod_5235 <- mkDebugOperation(mod_5235_inner, "mod_5235");
    Operation_IFC mod_5236_inner <- mkRepeatStatic(8);
    Operation_IFC mod_5236 <- mkDebugOperation(mod_5236_inner, "mod_5236");
    Operation_IFC mod_5237_inner <- mkFlatten(1);
    Operation_IFC mod_5237 <- mkDebugOperation(mod_5237_inner, "mod_5237");
    Operation_IFC mod_5238_inner <- mkFlatten(0);
    Operation_IFC mod_5238 <- mkDebugOperation(mod_5238_inner, "mod_5238");
    PMU_IFC mod_5239_bufferize <- mkPMU(1);
    Operation_IFC mod_5239_inner = mod_5239_bufferize.operation;
    Operation_IFC mod_5239 <- mkDebugOperation(mod_5239_inner, "mod_5239");
    Operation_IFC mod_5240_inner <- mkRepeatStatic(16);
    Operation_IFC mod_5240 <- mkDebugOperation(mod_5240_inner, "mod_5240");
    PMU_IFC mod_5241_bufferize <- mkPMU(2);
    Operation_IFC mod_5241_inner = mod_5241_bufferize.operation;
    Operation_IFC mod_5241 <- mkDebugOperation(mod_5241_inner, "mod_5241");
    Operation_IFC mod_5242_inner <- mkRepeatStatic(8);
    Operation_IFC mod_5242 <- mkDebugOperation(mod_5242_inner, "mod_5242");
    Operation_IFC mod_5243_inner <- mkFlatten(1);
    Operation_IFC mod_5243 <- mkDebugOperation(mod_5243_inner, "mod_5243");
    Operation_IFC mod_5244_inner <- mkFlatten(0);
    Operation_IFC mod_5244 <- mkDebugOperation(mod_5244_inner, "mod_5244");
    Operation_IFC mod_5245_inner <- mkRepeatStatic(16);
    Operation_IFC mod_5245 <- mkDebugOperation(mod_5245_inner, "mod_5245");
    Operation_IFC mod_5246_inner <- mkRepeatStatic(2);
    Operation_IFC mod_5246 <- mkDebugOperation(mod_5246_inner, "mod_5246");
    PMU_IFC mod_5247_bufferize <- mkPMU(2);
    Operation_IFC mod_5247_inner = mod_5247_bufferize.operation;
    Operation_IFC mod_5247 <- mkDebugOperation(mod_5247_inner, "mod_5247");
    rule rule_6732;
        ChannelMessage t;
        t <- mod_5230.get(0);
        mod_5229.put(0, t);
    endrule
    rule rule_6733;
        ChannelMessage t;
        t <- mod_5243.get(0);
        mod_5241.put(0, t);
    endrule
    rule rule_6734;
        ChannelMessage t;
        t <- mod_5238.get(0);
        mod_5237.put(0, t);
    endrule
    rule rule_6735;
        ChannelMessage t;
        t <- mod_5223.get(0);
        mod_5225.put(0, t);
    endrule
    rule rule_6736;
        ChannelMessage t;
        t <- mod_5212.get(3);
        mod_5213.put(0, t);
    endrule
    rule rule_6737;
        ChannelMessage t;
        t <- mod_5222.get(0);
        mod_5226.put(0, t);
    endrule
    rule rule_6738;
        ChannelMessage t;
        t <- mod_5213.get(1);
        mod_5214.put(0, t);
    endrule
    rule rule_6739;
        ChannelMessage t;
        t <- mod_5244.get(0);
        mod_5243.put(0, t);
    endrule
    rule rule_6740;
        ChannelMessage t;
        t <- mod_5211.get(0);
        mod_5247.put(0, t);
    endrule
    rule rule_6741;
        ChannelMessage t;
        t <- mod_5209.get(0);
        mod_5210.put(0, t);
    endrule
    rule rule_6742;
        ChannelMessage t;
        t <- mod_5211.get(1);
        mod_5212.put(0, t);
    endrule
    rule rule_6743;
        ChannelMessage t;
        t <- mod_5235.get(1);
        mod_5234.put(1, t);
    endrule
    rule rule_6744;
        ChannelMessage t;
        t <- mod_5241.get(0);
        mod_5242.put(0, t);
    endrule
    rule rule_6745;
        ChannelMessage t;
        t <- mod_5222.get(1);
        mod_5223.put(0, t);
    endrule
    rule rule_6746;
        ChannelMessage t;
        t <- mod_5231.get(0);
        mod_5219.put(1, t);
    endrule
    rule rule_6747;
        ChannelMessage t;
        t <- mod_5247.get(1);
        mod_5211.put(1, t);
    endrule
    rule rule_6748;
        ChannelMessage t;
        t <- mod_5239.get(0);
        mod_5240.put(0, t);
    endrule
    rule rule_6749;
        ChannelMessage t;
        t <- mod_5236.get(0);
        mod_5235.put(1, t);
    endrule
    rule rule_6750;
        ChannelMessage t;
        t <- mod_5240.get(0);
        mod_5239.put(1, t);
    endrule
    rule rule_6751;
        ChannelMessage t;
        t <- mod_5233.get(0);
        mod_5232.put(0, t);
    endrule
    rule rule_6752;
        ChannelMessage t;
        t <- mod_5225.get(0);
        mod_5225.put(1, t);
    endrule
    rule rule_6753;
        ChannelMessage t;
        t <- mod_5213.get(0);
        mod_5246.put(0, t);
    endrule
    rule rule_6754;
        ChannelMessage t;
        t <- mod_5223.get(1);
        mod_5224.put(1, t);
    endrule
    rule rule_6755;
        ChannelMessage t;
        t <- mod_5215.get(1);
        mod_5216.put(0, t);
    endrule
    rule rule_6756;
        ChannelMessage t;
        t <- mod_5210.get(0);
        mod_5211.put(0, t);
    endrule
    rule rule_6757;
        ChannelMessage t;
        t <- mod_5219.get(1);
        mod_5220.put(0, t);
    endrule
    rule rule_6758;
        ChannelMessage t;
        t <- mod_5246.get(0);
        mod_5213.put(1, t);
    endrule
    rule rule_6759;
        ChannelMessage t;
        t <- mod_5239.get(1);
        mod_5234.put(0, t);
    endrule
    rule rule_6760;
        ChannelMessage t;
        t <- mod_5225.get(1);
        mod_5223.put(1, t);
    endrule
    rule rule_6761;
        ChannelMessage t;
        t <- mod_5218.get(0);
        mod_5219.put(0, t);
    endrule
    rule rule_6762;
        ChannelMessage t;
        t <- mod_5214.get(0);
        mod_5239.put(0, t);
    endrule
    rule rule_6763;
        ChannelMessage t;
        t <- mod_5215.get(0);
        mod_5245.put(0, t);
    endrule
    rule rule_6764;
        ChannelMessage t;
        t <- mod_5234.get(0);
        mod_5233.put(0, t);
    endrule
    rule rule_6765;
        ChannelMessage t;
        t <- mod_5229.get(0);
        mod_5227.put(0, t);
    endrule
    rule rule_6766;
        ChannelMessage t;
        t <- mod_5214.get(1);
        mod_5215.put(0, t);
    endrule
    rule rule_6767;
        ChannelMessage t;
        t <- mod_5235.get(0);
        mod_5236.put(0, t);
    endrule
    rule rule_6768;
        ChannelMessage t;
        t <- mod_5227.get(1);
        mod_5220.put(1, t);
    endrule
    rule rule_6769;
        ChannelMessage t;
        t <- mod_5245.get(0);
        mod_5215.put(1, t);
    endrule
    rule rule_6770;
        ChannelMessage t;
        t <- mod_5226.get(1);
        mod_5222.put(1, t);
    endrule
    rule rule_6771;
        ChannelMessage t;
        t <- mod_5208.get(0);
        mod_5209.put(0, t);
    endrule
    rule rule_6772;
        ChannelMessage t;
        t <- mod_5216.get(0);
        mod_5217.put(0, t);
    endrule
    rule rule_6773;
        ChannelMessage t;
        t <- mod_5227.get(0);
        mod_5228.put(0, t);
    endrule
    rule rule_6774;
        ChannelMessage t;
        t <- mod_5237.get(0);
        mod_5235.put(0, t);
    endrule
    rule rule_6775;
        ChannelMessage t;
        t <- mod_5232.get(0);
        mod_5218.put(1, t);
    endrule
    rule rule_6776;
        ChannelMessage t;
        t <- mod_5217.get(0);
        mod_5218.put(0, t);
    endrule
    rule rule_6777;
        ChannelMessage t;
        t <- mod_5220.get(0);
        mod_5221.put(0, t);
    endrule
    rule rule_6778;
        ChannelMessage t;
        t <- mod_5247.get(0);
        mod_5247.put(1, t);
    endrule
    rule rule_6779;
        ChannelMessage t;
        t <- mod_5228.get(0);
        mod_5227.put(1, t);
    endrule
    rule rule_6780;
        ChannelMessage t;
        t <- mod_5219.get(0);
        mod_5231.put(0, t);
    endrule
    rule rule_6781;
        ChannelMessage t;
        t <- mod_5221.get(0);
        mod_5222.put(0, t);
    endrule
    rule rule_6782;
        ChannelMessage t;
        t <- mod_5241.get(1);
        mod_5216.put(1, t);
    endrule
    rule rule_6783;
        ChannelMessage t;
        t <- mod_5242.get(0);
        mod_5241.put(1, t);
    endrule
    rule rule_6784;
        ChannelMessage t;
        t <- mod_5226.get(0);
        mod_5226.put(1, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_5208.put(0, t);
        end
        if (i == 1) begin
            mod_5224.put(0, t);
        end
        if (i == 2) begin
            mod_5230.put(0, t);
        end
        if (i == 3) begin
            mod_5238.put(0, t);
        end
        if (i == 4) begin
            mod_5244.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_5212.get(0);
        end
        if (i == 3) begin
            t <- mod_5212.get(1);
        end
        if (i == 2) begin
            t <- mod_5212.get(2);
        end
        if (i == 1) begin
            t <- mod_5224.get(0);
        end

        return t;
    endmethod
endmodule

module mkStep(Empty);
    RamulatorArbiter_IFC#(0) ramulator_arbiter <- mkRamulatorArbiter(0);
    Operation_IFC mod_0_inner <- mkHypernode_6034;
    Operation_IFC mod_0 <- mkDebugOperation(mod_0_inner, "mod_0");
    Operation_IFC mod_41_inner <- mkHypernode_6035;
    Operation_IFC mod_41 <- mkDebugOperation(mod_41_inner, "mod_41");
    Operation_IFC mod_82_inner <- mkHypernode_6036;
    Operation_IFC mod_82 <- mkDebugOperation(mod_82_inner, "mod_82");
    Operation_IFC mod_123_inner <- mkHypernode_6037;
    Operation_IFC mod_123 <- mkDebugOperation(mod_123_inner, "mod_123");
    Operation_IFC mod_164_inner <- mkHypernode_6038;
    Operation_IFC mod_164 <- mkDebugOperation(mod_164_inner, "mod_164");
    Operation_IFC mod_205_inner <- mkHypernode_6039;
    Operation_IFC mod_205 <- mkDebugOperation(mod_205_inner, "mod_205");
    Operation_IFC mod_246_inner <- mkHypernode_6040;
    Operation_IFC mod_246 <- mkDebugOperation(mod_246_inner, "mod_246");
    Operation_IFC mod_287_inner <- mkHypernode_6041;
    Operation_IFC mod_287 <- mkDebugOperation(mod_287_inner, "mod_287");
    Operation_IFC mod_328_inner <- mkHypernode_6042;
    Operation_IFC mod_328 <- mkDebugOperation(mod_328_inner, "mod_328");
    Operation_IFC mod_369_inner <- mkHypernode_6043;
    Operation_IFC mod_369 <- mkDebugOperation(mod_369_inner, "mod_369");
    Operation_IFC mod_410_inner <- mkHypernode_6044;
    Operation_IFC mod_410 <- mkDebugOperation(mod_410_inner, "mod_410");
    Operation_IFC mod_451_inner <- mkHypernode_6045;
    Operation_IFC mod_451 <- mkDebugOperation(mod_451_inner, "mod_451");
    Operation_IFC mod_492_inner <- mkHypernode_6046;
    Operation_IFC mod_492 <- mkDebugOperation(mod_492_inner, "mod_492");
    Operation_IFC mod_533_inner <- mkHypernode_6047;
    Operation_IFC mod_533 <- mkDebugOperation(mod_533_inner, "mod_533");
    Operation_IFC mod_574_inner <- mkHypernode_6048;
    Operation_IFC mod_574 <- mkDebugOperation(mod_574_inner, "mod_574");
    Operation_IFC mod_615_inner <- mkHypernode_6049;
    Operation_IFC mod_615 <- mkDebugOperation(mod_615_inner, "mod_615");
    Operation_IFC mod_656_inner <- mkHypernode_6050;
    Operation_IFC mod_656 <- mkDebugOperation(mod_656_inner, "mod_656");
    Operation_IFC mod_697_inner <- mkHypernode_6051;
    Operation_IFC mod_697 <- mkDebugOperation(mod_697_inner, "mod_697");
    Operation_IFC mod_738_inner <- mkHypernode_6052;
    Operation_IFC mod_738 <- mkDebugOperation(mod_738_inner, "mod_738");
    Operation_IFC mod_779_inner <- mkHypernode_6053;
    Operation_IFC mod_779 <- mkDebugOperation(mod_779_inner, "mod_779");
    Operation_IFC mod_820_inner <- mkHypernode_6054;
    Operation_IFC mod_820 <- mkDebugOperation(mod_820_inner, "mod_820");
    Operation_IFC mod_861_inner <- mkHypernode_6055;
    Operation_IFC mod_861 <- mkDebugOperation(mod_861_inner, "mod_861");
    Operation_IFC mod_902_inner <- mkHypernode_6056;
    Operation_IFC mod_902 <- mkDebugOperation(mod_902_inner, "mod_902");
    Operation_IFC mod_943_inner <- mkHypernode_6057;
    Operation_IFC mod_943 <- mkDebugOperation(mod_943_inner, "mod_943");
    Operation_IFC mod_984_inner <- mkHypernode_6058;
    Operation_IFC mod_984 <- mkDebugOperation(mod_984_inner, "mod_984");
    Operation_IFC mod_1025_inner <- mkHypernode_6059;
    Operation_IFC mod_1025 <- mkDebugOperation(mod_1025_inner, "mod_1025");
    Operation_IFC mod_1066_inner <- mkHypernode_6060;
    Operation_IFC mod_1066 <- mkDebugOperation(mod_1066_inner, "mod_1066");
    Operation_IFC mod_1107_inner <- mkHypernode_6061;
    Operation_IFC mod_1107 <- mkDebugOperation(mod_1107_inner, "mod_1107");
    Operation_IFC mod_1148_inner <- mkHypernode_6062;
    Operation_IFC mod_1148 <- mkDebugOperation(mod_1148_inner, "mod_1148");
    Operation_IFC mod_1189_inner <- mkHypernode_6063;
    Operation_IFC mod_1189 <- mkDebugOperation(mod_1189_inner, "mod_1189");
    Operation_IFC mod_1230_inner <- mkHypernode_6064;
    Operation_IFC mod_1230 <- mkDebugOperation(mod_1230_inner, "mod_1230");
    Operation_IFC mod_1271_inner <- mkHypernode_6065;
    Operation_IFC mod_1271 <- mkDebugOperation(mod_1271_inner, "mod_1271");
    Operation_IFC mod_1312_inner <- mkHypernode_6066;
    Operation_IFC mod_1312 <- mkDebugOperation(mod_1312_inner, "mod_1312");
    Operation_IFC mod_1353_inner <- mkHypernode_6067;
    Operation_IFC mod_1353 <- mkDebugOperation(mod_1353_inner, "mod_1353");
    Operation_IFC mod_1394_inner <- mkHypernode_6068;
    Operation_IFC mod_1394 <- mkDebugOperation(mod_1394_inner, "mod_1394");
    Operation_IFC mod_1435_inner <- mkHypernode_6069;
    Operation_IFC mod_1435 <- mkDebugOperation(mod_1435_inner, "mod_1435");
    Operation_IFC mod_1476_inner <- mkHypernode_6070;
    Operation_IFC mod_1476 <- mkDebugOperation(mod_1476_inner, "mod_1476");
    Operation_IFC mod_1517_inner <- mkHypernode_6071;
    Operation_IFC mod_1517 <- mkDebugOperation(mod_1517_inner, "mod_1517");
    Operation_IFC mod_1558_inner <- mkHypernode_6072;
    Operation_IFC mod_1558 <- mkDebugOperation(mod_1558_inner, "mod_1558");
    Operation_IFC mod_1599_inner <- mkHypernode_6073;
    Operation_IFC mod_1599 <- mkDebugOperation(mod_1599_inner, "mod_1599");
    Operation_IFC mod_1640_inner <- mkHypernode_6074;
    Operation_IFC mod_1640 <- mkDebugOperation(mod_1640_inner, "mod_1640");
    Operation_IFC mod_1681_inner <- mkHypernode_6075;
    Operation_IFC mod_1681 <- mkDebugOperation(mod_1681_inner, "mod_1681");
    Operation_IFC mod_1722_inner <- mkHypernode_6076;
    Operation_IFC mod_1722 <- mkDebugOperation(mod_1722_inner, "mod_1722");
    Operation_IFC mod_1763_inner <- mkHypernode_6077;
    Operation_IFC mod_1763 <- mkDebugOperation(mod_1763_inner, "mod_1763");
    Operation_IFC mod_1804_inner <- mkHypernode_6078;
    Operation_IFC mod_1804 <- mkDebugOperation(mod_1804_inner, "mod_1804");
    Operation_IFC mod_1845_inner <- mkHypernode_6079;
    Operation_IFC mod_1845 <- mkDebugOperation(mod_1845_inner, "mod_1845");
    Operation_IFC mod_1886_inner <- mkHypernode_6080;
    Operation_IFC mod_1886 <- mkDebugOperation(mod_1886_inner, "mod_1886");
    Operation_IFC mod_1927_inner <- mkHypernode_6081;
    Operation_IFC mod_1927 <- mkDebugOperation(mod_1927_inner, "mod_1927");
    Operation_IFC mod_1968_inner <- mkHypernode_6082;
    Operation_IFC mod_1968 <- mkDebugOperation(mod_1968_inner, "mod_1968");
    Operation_IFC mod_2009_inner <- mkHypernode_6083;
    Operation_IFC mod_2009 <- mkDebugOperation(mod_2009_inner, "mod_2009");
    Operation_IFC mod_2050_inner <- mkHypernode_6084;
    Operation_IFC mod_2050 <- mkDebugOperation(mod_2050_inner, "mod_2050");
    Operation_IFC mod_2091_inner <- mkHypernode_6085;
    Operation_IFC mod_2091 <- mkDebugOperation(mod_2091_inner, "mod_2091");
    Operation_IFC mod_2132_inner <- mkHypernode_6086;
    Operation_IFC mod_2132 <- mkDebugOperation(mod_2132_inner, "mod_2132");
    Operation_IFC mod_2173_inner <- mkHypernode_6087;
    Operation_IFC mod_2173 <- mkDebugOperation(mod_2173_inner, "mod_2173");
    Operation_IFC mod_2214_inner <- mkHypernode_6088;
    Operation_IFC mod_2214 <- mkDebugOperation(mod_2214_inner, "mod_2214");
    Operation_IFC mod_2255_inner <- mkHypernode_6089;
    Operation_IFC mod_2255 <- mkDebugOperation(mod_2255_inner, "mod_2255");
    Operation_IFC mod_2296_inner <- mkHypernode_6090;
    Operation_IFC mod_2296 <- mkDebugOperation(mod_2296_inner, "mod_2296");
    Operation_IFC mod_2337_inner <- mkHypernode_6091;
    Operation_IFC mod_2337 <- mkDebugOperation(mod_2337_inner, "mod_2337");
    Operation_IFC mod_2378_inner <- mkHypernode_6092;
    Operation_IFC mod_2378 <- mkDebugOperation(mod_2378_inner, "mod_2378");
    Operation_IFC mod_2419_inner <- mkHypernode_6093;
    Operation_IFC mod_2419 <- mkDebugOperation(mod_2419_inner, "mod_2419");
    Operation_IFC mod_2460_inner <- mkHypernode_6094;
    Operation_IFC mod_2460 <- mkDebugOperation(mod_2460_inner, "mod_2460");
    Operation_IFC mod_2501_inner <- mkHypernode_6095;
    Operation_IFC mod_2501 <- mkDebugOperation(mod_2501_inner, "mod_2501");
    Operation_IFC mod_2542_inner <- mkHypernode_6096;
    Operation_IFC mod_2542 <- mkDebugOperation(mod_2542_inner, "mod_2542");
    Operation_IFC mod_2583_inner <- mkHypernode_6097;
    Operation_IFC mod_2583 <- mkDebugOperation(mod_2583_inner, "mod_2583");
    Operation_IFC mod_2624_inner <- mkHypernode_6098;
    Operation_IFC mod_2624 <- mkDebugOperation(mod_2624_inner, "mod_2624");
    Operation_IFC mod_2665_inner <- mkHypernode_6099;
    Operation_IFC mod_2665 <- mkDebugOperation(mod_2665_inner, "mod_2665");
    Operation_IFC mod_2706_inner <- mkHypernode_6100;
    Operation_IFC mod_2706 <- mkDebugOperation(mod_2706_inner, "mod_2706");
    Operation_IFC mod_2747_inner <- mkHypernode_6101;
    Operation_IFC mod_2747 <- mkDebugOperation(mod_2747_inner, "mod_2747");
    Operation_IFC mod_2788_inner <- mkHypernode_6102;
    Operation_IFC mod_2788 <- mkDebugOperation(mod_2788_inner, "mod_2788");
    Operation_IFC mod_2829_inner <- mkHypernode_6103;
    Operation_IFC mod_2829 <- mkDebugOperation(mod_2829_inner, "mod_2829");
    Operation_IFC mod_2870_inner <- mkHypernode_6104;
    Operation_IFC mod_2870 <- mkDebugOperation(mod_2870_inner, "mod_2870");
    Operation_IFC mod_2911_inner <- mkHypernode_6105;
    Operation_IFC mod_2911 <- mkDebugOperation(mod_2911_inner, "mod_2911");
    Operation_IFC mod_2952_inner <- mkHypernode_6106;
    Operation_IFC mod_2952 <- mkDebugOperation(mod_2952_inner, "mod_2952");
    Operation_IFC mod_2993_inner <- mkHypernode_6107;
    Operation_IFC mod_2993 <- mkDebugOperation(mod_2993_inner, "mod_2993");
    Operation_IFC mod_3034_inner <- mkHypernode_6108;
    Operation_IFC mod_3034 <- mkDebugOperation(mod_3034_inner, "mod_3034");
    Operation_IFC mod_3075_inner <- mkHypernode_6109;
    Operation_IFC mod_3075 <- mkDebugOperation(mod_3075_inner, "mod_3075");
    Operation_IFC mod_3116_inner <- mkHypernode_6110;
    Operation_IFC mod_3116 <- mkDebugOperation(mod_3116_inner, "mod_3116");
    Operation_IFC mod_3157_inner <- mkHypernode_6111;
    Operation_IFC mod_3157 <- mkDebugOperation(mod_3157_inner, "mod_3157");
    Operation_IFC mod_3198_inner <- mkHypernode_6112;
    Operation_IFC mod_3198 <- mkDebugOperation(mod_3198_inner, "mod_3198");
    Operation_IFC mod_3239_inner <- mkHypernode_6113;
    Operation_IFC mod_3239 <- mkDebugOperation(mod_3239_inner, "mod_3239");
    Operation_IFC mod_3280_inner <- mkHypernode_6114;
    Operation_IFC mod_3280 <- mkDebugOperation(mod_3280_inner, "mod_3280");
    Operation_IFC mod_3321_inner <- mkHypernode_6115;
    Operation_IFC mod_3321 <- mkDebugOperation(mod_3321_inner, "mod_3321");
    Operation_IFC mod_3362_inner <- mkHypernode_6116;
    Operation_IFC mod_3362 <- mkDebugOperation(mod_3362_inner, "mod_3362");
    Operation_IFC mod_3403_inner <- mkHypernode_6117;
    Operation_IFC mod_3403 <- mkDebugOperation(mod_3403_inner, "mod_3403");
    Operation_IFC mod_3444_inner <- mkHypernode_6118;
    Operation_IFC mod_3444 <- mkDebugOperation(mod_3444_inner, "mod_3444");
    Operation_IFC mod_3485_inner <- mkHypernode_6119;
    Operation_IFC mod_3485 <- mkDebugOperation(mod_3485_inner, "mod_3485");
    Operation_IFC mod_3526_inner <- mkHypernode_6120;
    Operation_IFC mod_3526 <- mkDebugOperation(mod_3526_inner, "mod_3526");
    Operation_IFC mod_3567_inner <- mkHypernode_6121;
    Operation_IFC mod_3567 <- mkDebugOperation(mod_3567_inner, "mod_3567");
    Operation_IFC mod_3608_inner <- mkHypernode_6122;
    Operation_IFC mod_3608 <- mkDebugOperation(mod_3608_inner, "mod_3608");
    Operation_IFC mod_3649_inner <- mkHypernode_6123;
    Operation_IFC mod_3649 <- mkDebugOperation(mod_3649_inner, "mod_3649");
    Operation_IFC mod_3690_inner <- mkHypernode_6124;
    Operation_IFC mod_3690 <- mkDebugOperation(mod_3690_inner, "mod_3690");
    Operation_IFC mod_3731_inner <- mkHypernode_6125;
    Operation_IFC mod_3731 <- mkDebugOperation(mod_3731_inner, "mod_3731");
    Operation_IFC mod_3772_inner <- mkHypernode_6126;
    Operation_IFC mod_3772 <- mkDebugOperation(mod_3772_inner, "mod_3772");
    Operation_IFC mod_3813_inner <- mkHypernode_6127;
    Operation_IFC mod_3813 <- mkDebugOperation(mod_3813_inner, "mod_3813");
    Operation_IFC mod_3854_inner <- mkHypernode_6128;
    Operation_IFC mod_3854 <- mkDebugOperation(mod_3854_inner, "mod_3854");
    Operation_IFC mod_3895_inner <- mkHypernode_6129;
    Operation_IFC mod_3895 <- mkDebugOperation(mod_3895_inner, "mod_3895");
    Operation_IFC mod_3936_inner <- mkHypernode_6130;
    Operation_IFC mod_3936 <- mkDebugOperation(mod_3936_inner, "mod_3936");
    Operation_IFC mod_3977_inner <- mkHypernode_6131;
    Operation_IFC mod_3977 <- mkDebugOperation(mod_3977_inner, "mod_3977");
    Operation_IFC mod_4018_inner <- mkHypernode_6132;
    Operation_IFC mod_4018 <- mkDebugOperation(mod_4018_inner, "mod_4018");
    Operation_IFC mod_4059_inner <- mkHypernode_6133;
    Operation_IFC mod_4059 <- mkDebugOperation(mod_4059_inner, "mod_4059");
    Operation_IFC mod_4100_inner <- mkHypernode_6134;
    Operation_IFC mod_4100 <- mkDebugOperation(mod_4100_inner, "mod_4100");
    Operation_IFC mod_4141_inner <- mkHypernode_6135;
    Operation_IFC mod_4141 <- mkDebugOperation(mod_4141_inner, "mod_4141");
    Operation_IFC mod_4182_inner <- mkHypernode_6136;
    Operation_IFC mod_4182 <- mkDebugOperation(mod_4182_inner, "mod_4182");
    Operation_IFC mod_4223_inner <- mkHypernode_6137;
    Operation_IFC mod_4223 <- mkDebugOperation(mod_4223_inner, "mod_4223");
    Operation_IFC mod_4264_inner <- mkHypernode_6138;
    Operation_IFC mod_4264 <- mkDebugOperation(mod_4264_inner, "mod_4264");
    Operation_IFC mod_4305_inner <- mkHypernode_6139;
    Operation_IFC mod_4305 <- mkDebugOperation(mod_4305_inner, "mod_4305");
    Operation_IFC mod_4346_inner <- mkHypernode_6140;
    Operation_IFC mod_4346 <- mkDebugOperation(mod_4346_inner, "mod_4346");
    Operation_IFC mod_4387_inner <- mkHypernode_6141;
    Operation_IFC mod_4387 <- mkDebugOperation(mod_4387_inner, "mod_4387");
    Operation_IFC mod_4428_inner <- mkHypernode_6142;
    Operation_IFC mod_4428 <- mkDebugOperation(mod_4428_inner, "mod_4428");
    Operation_IFC mod_4469_inner <- mkHypernode_6143;
    Operation_IFC mod_4469 <- mkDebugOperation(mod_4469_inner, "mod_4469");
    Operation_IFC mod_4510_inner <- mkHypernode_6144;
    Operation_IFC mod_4510 <- mkDebugOperation(mod_4510_inner, "mod_4510");
    Operation_IFC mod_4551_inner <- mkHypernode_6145;
    Operation_IFC mod_4551 <- mkDebugOperation(mod_4551_inner, "mod_4551");
    Operation_IFC mod_4592_inner <- mkHypernode_6146;
    Operation_IFC mod_4592 <- mkDebugOperation(mod_4592_inner, "mod_4592");
    Operation_IFC mod_4633_inner <- mkHypernode_6147;
    Operation_IFC mod_4633 <- mkDebugOperation(mod_4633_inner, "mod_4633");
    Operation_IFC mod_4674_inner <- mkHypernode_6148;
    Operation_IFC mod_4674 <- mkDebugOperation(mod_4674_inner, "mod_4674");
    Operation_IFC mod_4715_inner <- mkHypernode_6149;
    Operation_IFC mod_4715 <- mkDebugOperation(mod_4715_inner, "mod_4715");
    Operation_IFC mod_4756_inner <- mkHypernode_6150;
    Operation_IFC mod_4756 <- mkDebugOperation(mod_4756_inner, "mod_4756");
    Operation_IFC mod_4797_inner <- mkHypernode_6151;
    Operation_IFC mod_4797 <- mkDebugOperation(mod_4797_inner, "mod_4797");
    Operation_IFC mod_4838_inner <- mkHypernode_6152;
    Operation_IFC mod_4838 <- mkDebugOperation(mod_4838_inner, "mod_4838");
    Operation_IFC mod_4879_inner <- mkHypernode_6153;
    Operation_IFC mod_4879 <- mkDebugOperation(mod_4879_inner, "mod_4879");
    Operation_IFC mod_4920_inner <- mkHypernode_6154;
    Operation_IFC mod_4920 <- mkDebugOperation(mod_4920_inner, "mod_4920");
    Operation_IFC mod_4961_inner <- mkHypernode_6155;
    Operation_IFC mod_4961 <- mkDebugOperation(mod_4961_inner, "mod_4961");
    Operation_IFC mod_5002_inner <- mkHypernode_6156;
    Operation_IFC mod_5002 <- mkDebugOperation(mod_5002_inner, "mod_5002");
    Operation_IFC mod_5043_inner <- mkHypernode_6157;
    Operation_IFC mod_5043 <- mkDebugOperation(mod_5043_inner, "mod_5043");
    Operation_IFC mod_5084_inner <- mkHypernode_6158;
    Operation_IFC mod_5084 <- mkDebugOperation(mod_5084_inner, "mod_5084");
    Operation_IFC mod_5125_inner <- mkHypernode_6159;
    Operation_IFC mod_5125 <- mkDebugOperation(mod_5125_inner, "mod_5125");
    Operation_IFC mod_5166_inner <- mkHypernode_6160;
    Operation_IFC mod_5166 <- mkDebugOperation(mod_5166_inner, "mod_5166");
    Operation_IFC mod_5207_inner <- mkHypernode_6161;
    Operation_IFC mod_5207 <- mkDebugOperation(mod_5207_inner, "mod_5207");
    Operation_IFC mod_5248_inner <- mkFlatten(0);
    Operation_IFC mod_5248 <- mkDebugOperation(mod_5248_inner, "mod_5248");
    Operation_IFC mod_5249_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5249 <- mkDebugOperation(mod_5249_inner, "mod_5249");
    Operation_IFC mod_5250_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5250 <- mkDebugOperation(mod_5250_inner, "mod_5250");
    Operation_IFC mod_5251_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5251 <- mkDebugOperation(mod_5251_inner, "mod_5251");
    Operation_IFC mod_5252_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5252 <- mkDebugOperation(mod_5252_inner, "mod_5252");
    Operation_IFC mod_5253_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5253 <- mkDebugOperation(mod_5253_inner, "mod_5253");
    Operation_IFC mod_5254_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5254 <- mkDebugOperation(mod_5254_inner, "mod_5254");
    Operation_IFC mod_5255_inner <- mkPrinter("mod_5255");
    Operation_IFC mod_5255 <- mkDebugOperation(mod_5255_inner, "mod_5255");
    Operation_IFC mod_5256_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5256 <- mkDebugOperation(mod_5256_inner, "mod_5256");
    Operation_IFC mod_5257_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5257 <- mkDebugOperation(mod_5257_inner, "mod_5257");
    Operation_IFC mod_5258_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5258 <- mkDebugOperation(mod_5258_inner, "mod_5258");
    Operation_IFC mod_5259_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5259 <- mkDebugOperation(mod_5259_inner, "mod_5259");
    Operation_IFC mod_5260_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5260 <- mkDebugOperation(mod_5260_inner, "mod_5260");
    Operation_IFC mod_5261_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5261 <- mkDebugOperation(mod_5261_inner, "mod_5261");
    Operation_IFC mod_5262_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5262 <- mkDebugOperation(mod_5262_inner, "mod_5262");
    Operation_IFC mod_5263_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5263 <- mkDebugOperation(mod_5263_inner, "mod_5263");
    Operation_IFC mod_5264_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5264 <- mkDebugOperation(mod_5264_inner, "mod_5264");
    Operation_IFC mod_5265_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5265 <- mkDebugOperation(mod_5265_inner, "mod_5265");
    Operation_IFC mod_5266_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5266 <- mkDebugOperation(mod_5266_inner, "mod_5266");
    Operation_IFC mod_5267_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5267 <- mkDebugOperation(mod_5267_inner, "mod_5267");
    Operation_IFC mod_5268_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5268 <- mkDebugOperation(mod_5268_inner, "mod_5268");
    Operation_IFC mod_5269_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5269 <- mkDebugOperation(mod_5269_inner, "mod_5269");
    Operation_IFC mod_5270_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5270 <- mkDebugOperation(mod_5270_inner, "mod_5270");
    Operation_IFC mod_5271_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5271 <- mkDebugOperation(mod_5271_inner, "mod_5271");
    Operation_IFC mod_5272_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5272 <- mkDebugOperation(mod_5272_inner, "mod_5272");
    Operation_IFC mod_5273_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5273 <- mkDebugOperation(mod_5273_inner, "mod_5273");
    Operation_IFC mod_5274_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5274 <- mkDebugOperation(mod_5274_inner, "mod_5274");
    Operation_IFC mod_5275_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5275 <- mkDebugOperation(mod_5275_inner, "mod_5275");
    Operation_IFC mod_5276_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5276 <- mkDebugOperation(mod_5276_inner, "mod_5276");
    Operation_IFC mod_5277_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5277 <- mkDebugOperation(mod_5277_inner, "mod_5277");
    Operation_IFC mod_5278_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5278 <- mkDebugOperation(mod_5278_inner, "mod_5278");
    Operation_IFC mod_5279_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5279 <- mkDebugOperation(mod_5279_inner, "mod_5279");
    Operation_IFC mod_5280_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5280 <- mkDebugOperation(mod_5280_inner, "mod_5280");
    Operation_IFC mod_5281_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5281 <- mkDebugOperation(mod_5281_inner, "mod_5281");
    Operation_IFC mod_5282_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5282 <- mkDebugOperation(mod_5282_inner, "mod_5282");
    Operation_IFC mod_5283_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5283 <- mkDebugOperation(mod_5283_inner, "mod_5283");
    Operation_IFC mod_5284_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5284 <- mkDebugOperation(mod_5284_inner, "mod_5284");
    Operation_IFC mod_5285_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5285 <- mkDebugOperation(mod_5285_inner, "mod_5285");
    Operation_IFC mod_5286_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5286 <- mkDebugOperation(mod_5286_inner, "mod_5286");
    Operation_IFC mod_5287_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5287 <- mkDebugOperation(mod_5287_inner, "mod_5287");
    Operation_IFC mod_5288_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5288 <- mkDebugOperation(mod_5288_inner, "mod_5288");
    Operation_IFC mod_5289_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5289 <- mkDebugOperation(mod_5289_inner, "mod_5289");
    Operation_IFC mod_5290_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5290 <- mkDebugOperation(mod_5290_inner, "mod_5290");
    Operation_IFC mod_5291_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5291 <- mkDebugOperation(mod_5291_inner, "mod_5291");
    Operation_IFC mod_5292_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5292 <- mkDebugOperation(mod_5292_inner, "mod_5292");
    Operation_IFC mod_5293_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5293 <- mkDebugOperation(mod_5293_inner, "mod_5293");
    Operation_IFC mod_5294_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5294 <- mkDebugOperation(mod_5294_inner, "mod_5294");
    Operation_IFC mod_5295_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5295 <- mkDebugOperation(mod_5295_inner, "mod_5295");
    Operation_IFC mod_5296_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5296 <- mkDebugOperation(mod_5296_inner, "mod_5296");
    Operation_IFC mod_5297_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5297 <- mkDebugOperation(mod_5297_inner, "mod_5297");
    Operation_IFC mod_5298_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5298 <- mkDebugOperation(mod_5298_inner, "mod_5298");
    Operation_IFC mod_5299_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5299 <- mkDebugOperation(mod_5299_inner, "mod_5299");
    Operation_IFC mod_5300_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5300 <- mkDebugOperation(mod_5300_inner, "mod_5300");
    Operation_IFC mod_5301_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5301 <- mkDebugOperation(mod_5301_inner, "mod_5301");
    Operation_IFC mod_5302_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5302 <- mkDebugOperation(mod_5302_inner, "mod_5302");
    Operation_IFC mod_5303_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5303 <- mkDebugOperation(mod_5303_inner, "mod_5303");
    Operation_IFC mod_5304_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5304 <- mkDebugOperation(mod_5304_inner, "mod_5304");
    Operation_IFC mod_5305_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5305 <- mkDebugOperation(mod_5305_inner, "mod_5305");
    Operation_IFC mod_5306_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5306 <- mkDebugOperation(mod_5306_inner, "mod_5306");
    Operation_IFC mod_5307_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5307 <- mkDebugOperation(mod_5307_inner, "mod_5307");
    Operation_IFC mod_5308_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5308 <- mkDebugOperation(mod_5308_inner, "mod_5308");
    Partition_IFC#(128) mod_5309_inner <- mkPartition(0, 128);
    Operation_IFC mod_5309 <- mkDebugOperation(mod_5309_inner.op, "mod_5309");
    Operation_IFC mod_5310_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5310 <- mkDebugOperation(mod_5310_inner, "mod_5310");
    Operation_IFC mod_5311_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5311 <- mkDebugOperation(mod_5311_inner, "mod_5311");
    Operation_IFC mod_5312_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5312 <- mkDebugOperation(mod_5312_inner, "mod_5312");
    Reassemble_IFC#(128) mod_5313_inner <- mkReassemble(128);
    Operation_IFC mod_5313 <- mkDebugOperation(mod_5313_inner.op, "mod_5313");
    Operation_IFC mod_5314_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5314 <- mkDebugOperation(mod_5314_inner, "mod_5314");
    Operation_IFC mod_5315_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5315 <- mkDebugOperation(mod_5315_inner, "mod_5315");
    Operation_IFC mod_5316_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5316 <- mkDebugOperation(mod_5316_inner, "mod_5316");
    Operation_IFC mod_5317_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5317 <- mkDebugOperation(mod_5317_inner, "mod_5317");
    Operation_IFC mod_5318_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5318 <- mkDebugOperation(mod_5318_inner, "mod_5318");
    Operation_IFC mod_5319_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5319 <- mkDebugOperation(mod_5319_inner, "mod_5319");
    Operation_IFC mod_5320_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5320 <- mkDebugOperation(mod_5320_inner, "mod_5320");
    Operation_IFC mod_5321_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5321 <- mkDebugOperation(mod_5321_inner, "mod_5321");
    Operation_IFC mod_5322_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5322 <- mkDebugOperation(mod_5322_inner, "mod_5322");
    Operation_IFC mod_5323_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5323 <- mkDebugOperation(mod_5323_inner, "mod_5323");
    Operation_IFC mod_5324_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5324 <- mkDebugOperation(mod_5324_inner, "mod_5324");
    Operation_IFC mod_5325_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5325 <- mkDebugOperation(mod_5325_inner, "mod_5325");
    PMU_IFC mod_5326_bufferize <- mkPMU(2);
    Operation_IFC mod_5326_inner = mod_5326_bufferize.operation;
    Operation_IFC mod_5326 <- mkDebugOperation(mod_5326_inner, "mod_5326");
    Operation_IFC mod_5327_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5327 <- mkDebugOperation(mod_5327_inner, "mod_5327");
    Operation_IFC mod_5328_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5328 <- mkDebugOperation(mod_5328_inner, "mod_5328");
    Operation_IFC mod_5329_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5329 <- mkDebugOperation(mod_5329_inner, "mod_5329");
    Operation_IFC mod_5330_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5330 <- mkDebugOperation(mod_5330_inner, "mod_5330");
    Operation_IFC mod_5331_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5331 <- mkDebugOperation(mod_5331_inner, "mod_5331");
    Operation_IFC mod_5332_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5332 <- mkDebugOperation(mod_5332_inner, "mod_5332");
    Operation_IFC mod_5333_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5333 <- mkDebugOperation(mod_5333_inner, "mod_5333");
    Operation_IFC mod_5334_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5334 <- mkDebugOperation(mod_5334_inner, "mod_5334");
    Operation_IFC mod_5335_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5335 <- mkDebugOperation(mod_5335_inner, "mod_5335");
    Operation_IFC mod_5336_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5336 <- mkDebugOperation(mod_5336_inner, "mod_5336");
    Operation_IFC mod_5337_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5337 <- mkDebugOperation(mod_5337_inner, "mod_5337");
    Operation_IFC mod_5338_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5338 <- mkDebugOperation(mod_5338_inner, "mod_5338");
    Operation_IFC mod_5339_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5339 <- mkDebugOperation(mod_5339_inner, "mod_5339");
    Operation_IFC mod_5340_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5340 <- mkDebugOperation(mod_5340_inner, "mod_5340");
    Operation_IFC mod_5341_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5341 <- mkDebugOperation(mod_5341_inner, "mod_5341");
    Operation_IFC mod_5342_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5342 <- mkDebugOperation(mod_5342_inner, "mod_5342");
    Operation_IFC mod_5343_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5343 <- mkDebugOperation(mod_5343_inner, "mod_5343");
    Operation_IFC mod_5344_inner <- mkRandomOffChipLoad(Cons(64, Cons(1, Cons(1, Cons(1, Cons(1, Cons(1, Nil)))))));
    Operation_IFC mod_5344 <- mkDebugOperation(mod_5344_inner, "mod_5344");
    Operation_IFC mod_5345_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5345 <- mkDebugOperation(mod_5345_inner, "mod_5345");
    Operation_IFC mod_5346_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5346 <- mkDebugOperation(mod_5346_inner, "mod_5346");
    Operation_IFC mod_5347_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5347 <- mkDebugOperation(mod_5347_inner, "mod_5347");
    Operation_IFC mod_5348_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5348 <- mkDebugOperation(mod_5348_inner, "mod_5348");
    Operation_IFC mod_5349_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5349 <- mkDebugOperation(mod_5349_inner, "mod_5349");
    Operation_IFC mod_5350_inner <- mkRandomSelectGen;
    Operation_IFC mod_5350 <- mkDebugOperation(mod_5350_inner, "mod_5350");
    Operation_IFC mod_5351_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5351 <- mkDebugOperation(mod_5351_inner, "mod_5351");
    Operation_IFC mod_5352_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5352 <- mkDebugOperation(mod_5352_inner, "mod_5352");
    Operation_IFC mod_5353_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5353 <- mkDebugOperation(mod_5353_inner, "mod_5353");
    Operation_IFC mod_5354_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5354 <- mkDebugOperation(mod_5354_inner, "mod_5354");
    Operation_IFC mod_5355_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5355 <- mkDebugOperation(mod_5355_inner, "mod_5355");
    Operation_IFC mod_5356_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5356 <- mkDebugOperation(mod_5356_inner, "mod_5356");
    Operation_IFC mod_5357_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5357 <- mkDebugOperation(mod_5357_inner, "mod_5357");
    Operation_IFC mod_5358_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5358 <- mkDebugOperation(mod_5358_inner, "mod_5358");
    Operation_IFC mod_5359_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5359 <- mkDebugOperation(mod_5359_inner, "mod_5359");
    Operation_IFC mod_5360_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5360 <- mkDebugOperation(mod_5360_inner, "mod_5360");
    Operation_IFC mod_5361_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5361 <- mkDebugOperation(mod_5361_inner, "mod_5361");
    Operation_IFC mod_5362_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5362 <- mkDebugOperation(mod_5362_inner, "mod_5362");
    Operation_IFC mod_5363_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5363 <- mkDebugOperation(mod_5363_inner, "mod_5363");
    Operation_IFC mod_5364_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5364 <- mkDebugOperation(mod_5364_inner, "mod_5364");
    Operation_IFC mod_5365_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5365 <- mkDebugOperation(mod_5365_inner, "mod_5365");
    Operation_IFC mod_5366_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5366 <- mkDebugOperation(mod_5366_inner, "mod_5366");
    Operation_IFC mod_5367_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5367 <- mkDebugOperation(mod_5367_inner, "mod_5367");
    Operation_IFC mod_5368_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5368 <- mkDebugOperation(mod_5368_inner, "mod_5368");
    Operation_IFC mod_5369_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5369 <- mkDebugOperation(mod_5369_inner, "mod_5369");
    Operation_IFC mod_5370_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5370 <- mkDebugOperation(mod_5370_inner, "mod_5370");
    Operation_IFC mod_5371_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5371 <- mkDebugOperation(mod_5371_inner, "mod_5371");
    Operation_IFC mod_5372_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_5372 <- mkDebugOperation(mod_5372_inner, "mod_5372");
    Operation_IFC mod_5373_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5373 <- mkDebugOperation(mod_5373_inner, "mod_5373");
    Operation_IFC mod_5374_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5374 <- mkDebugOperation(mod_5374_inner, "mod_5374");
    Operation_IFC mod_5375_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5375 <- mkDebugOperation(mod_5375_inner, "mod_5375");
    Operation_IFC mod_5376_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5376 <- mkDebugOperation(mod_5376_inner, "mod_5376");
    Operation_IFC mod_5377_inner <- mkRepeatStatic(1);
    Operation_IFC mod_5377 <- mkDebugOperation(mod_5377_inner, "mod_5377");
    Operation_IFC mod_5378_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5378 <- mkDebugOperation(mod_5378_inner, "mod_5378");
    Operation_IFC mod_5379_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5379 <- mkDebugOperation(mod_5379_inner, "mod_5379");
    Operation_IFC mod_5380_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5380 <- mkDebugOperation(mod_5380_inner, "mod_5380");
    Operation_IFC mod_5381_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5381 <- mkDebugOperation(mod_5381_inner, "mod_5381");
    Operation_IFC mod_5382_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5382 <- mkDebugOperation(mod_5382_inner, "mod_5382");
    Operation_IFC mod_5383_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5383 <- mkDebugOperation(mod_5383_inner, "mod_5383");
    Operation_IFC mod_5384_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5384 <- mkDebugOperation(mod_5384_inner, "mod_5384");
    Operation_IFC mod_5385_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5385 <- mkDebugOperation(mod_5385_inner, "mod_5385");
    Operation_IFC mod_5386_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5386 <- mkDebugOperation(mod_5386_inner, "mod_5386");
    Operation_IFC mod_5387_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5387 <- mkDebugOperation(mod_5387_inner, "mod_5387");
    Operation_IFC mod_5388_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5388 <- mkDebugOperation(mod_5388_inner, "mod_5388");
    Operation_IFC mod_5389_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5389 <- mkDebugOperation(mod_5389_inner, "mod_5389");
    Operation_IFC mod_5390_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5390 <- mkDebugOperation(mod_5390_inner, "mod_5390");
    Operation_IFC mod_5391_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5391 <- mkDebugOperation(mod_5391_inner, "mod_5391");
    Operation_IFC mod_5392_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5392 <- mkDebugOperation(mod_5392_inner, "mod_5392");
    Operation_IFC mod_5393_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5393 <- mkDebugOperation(mod_5393_inner, "mod_5393");
    Operation_IFC mod_5394_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5394 <- mkDebugOperation(mod_5394_inner, "mod_5394");
    Operation_IFC mod_5395_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5395 <- mkDebugOperation(mod_5395_inner, "mod_5395");
    Operation_IFC mod_5396_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5396 <- mkDebugOperation(mod_5396_inner, "mod_5396");
    Operation_IFC mod_5397_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5397 <- mkDebugOperation(mod_5397_inner, "mod_5397");
    Operation_IFC mod_5398_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5398 <- mkDebugOperation(mod_5398_inner, "mod_5398");
    Operation_IFC mod_5399_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5399 <- mkDebugOperation(mod_5399_inner, "mod_5399");
    Operation_IFC mod_5400_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5400 <- mkDebugOperation(mod_5400_inner, "mod_5400");
    Operation_IFC mod_5401_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5401 <- mkDebugOperation(mod_5401_inner, "mod_5401");
    Operation_IFC mod_5402_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5402 <- mkDebugOperation(mod_5402_inner, "mod_5402");
    Operation_IFC mod_5403_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5403 <- mkDebugOperation(mod_5403_inner, "mod_5403");
    Operation_IFC mod_5404_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5404 <- mkDebugOperation(mod_5404_inner, "mod_5404");
    Operation_IFC mod_5405_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5405 <- mkDebugOperation(mod_5405_inner, "mod_5405");
    Operation_IFC mod_5406_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5406 <- mkDebugOperation(mod_5406_inner, "mod_5406");
    Operation_IFC mod_5407_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5407 <- mkDebugOperation(mod_5407_inner, "mod_5407");
    Operation_IFC mod_5408_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5408 <- mkDebugOperation(mod_5408_inner, "mod_5408");
    Operation_IFC mod_5409_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5409 <- mkDebugOperation(mod_5409_inner, "mod_5409");
    Operation_IFC mod_5410_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5410 <- mkDebugOperation(mod_5410_inner, "mod_5410");
    Operation_IFC mod_5411_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5411 <- mkDebugOperation(mod_5411_inner, "mod_5411");
    Operation_IFC mod_5412_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5412 <- mkDebugOperation(mod_5412_inner, "mod_5412");
    Operation_IFC mod_5413_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5413 <- mkDebugOperation(mod_5413_inner, "mod_5413");
    Operation_IFC mod_5414_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5414 <- mkDebugOperation(mod_5414_inner, "mod_5414");
    Operation_IFC mod_5415_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5415 <- mkDebugOperation(mod_5415_inner, "mod_5415");
    Operation_IFC mod_5416_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5416 <- mkDebugOperation(mod_5416_inner, "mod_5416");
    Operation_IFC mod_5417_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5417 <- mkDebugOperation(mod_5417_inner, "mod_5417");
    Operation_IFC mod_5418_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5418 <- mkDebugOperation(mod_5418_inner, "mod_5418");
    Operation_IFC mod_5419_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5419 <- mkDebugOperation(mod_5419_inner, "mod_5419");
    Operation_IFC mod_5420_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5420 <- mkDebugOperation(mod_5420_inner, "mod_5420");
    Operation_IFC mod_5421_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5421 <- mkDebugOperation(mod_5421_inner, "mod_5421");
    Operation_IFC mod_5422_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5422 <- mkDebugOperation(mod_5422_inner, "mod_5422");
    Operation_IFC mod_5423_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5423 <- mkDebugOperation(mod_5423_inner, "mod_5423");
    Operation_IFC mod_5424_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5424 <- mkDebugOperation(mod_5424_inner, "mod_5424");
    Operation_IFC mod_5425_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5425 <- mkDebugOperation(mod_5425_inner, "mod_5425");
    Operation_IFC mod_5426_inner <- mkRandomSelectGen;
    Operation_IFC mod_5426 <- mkDebugOperation(mod_5426_inner, "mod_5426");
    Operation_IFC mod_5427_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5427 <- mkDebugOperation(mod_5427_inner, "mod_5427");
    Operation_IFC mod_5428_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5428 <- mkDebugOperation(mod_5428_inner, "mod_5428");
    Operation_IFC mod_5429_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5429 <- mkDebugOperation(mod_5429_inner, "mod_5429");
    Operation_IFC mod_5430_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5430 <- mkDebugOperation(mod_5430_inner, "mod_5430");
    Operation_IFC mod_5431_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5431 <- mkDebugOperation(mod_5431_inner, "mod_5431");
    Operation_IFC mod_5432_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5432 <- mkDebugOperation(mod_5432_inner, "mod_5432");
    Operation_IFC mod_5433_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5433 <- mkDebugOperation(mod_5433_inner, "mod_5433");
    Operation_IFC mod_5434_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5434 <- mkDebugOperation(mod_5434_inner, "mod_5434");
    Operation_IFC mod_5435_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5435 <- mkDebugOperation(mod_5435_inner, "mod_5435");
    Operation_IFC mod_5436_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5436 <- mkDebugOperation(mod_5436_inner, "mod_5436");
    Operation_IFC mod_5437_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5437 <- mkDebugOperation(mod_5437_inner, "mod_5437");
    Operation_IFC mod_5438_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5438 <- mkDebugOperation(mod_5438_inner, "mod_5438");
    Operation_IFC mod_5439_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5439 <- mkDebugOperation(mod_5439_inner, "mod_5439");
    Operation_IFC mod_5440_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5440 <- mkDebugOperation(mod_5440_inner, "mod_5440");
    Operation_IFC mod_5441_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5441 <- mkDebugOperation(mod_5441_inner, "mod_5441");
    Operation_IFC mod_5442_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5442 <- mkDebugOperation(mod_5442_inner, "mod_5442");
    Operation_IFC mod_5443_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5443 <- mkDebugOperation(mod_5443_inner, "mod_5443");
    Operation_IFC mod_5444_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5444 <- mkDebugOperation(mod_5444_inner, "mod_5444");
    Operation_IFC mod_5445_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5445 <- mkDebugOperation(mod_5445_inner, "mod_5445");
    Operation_IFC mod_5446_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5446 <- mkDebugOperation(mod_5446_inner, "mod_5446");
    Operation_IFC mod_5447_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5447 <- mkDebugOperation(mod_5447_inner, "mod_5447");
    Operation_IFC mod_5448_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5448 <- mkDebugOperation(mod_5448_inner, "mod_5448");
    Operation_IFC mod_5449_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5449 <- mkDebugOperation(mod_5449_inner, "mod_5449");
    Operation_IFC mod_5450_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5450 <- mkDebugOperation(mod_5450_inner, "mod_5450");
    Operation_IFC mod_5451_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5451 <- mkDebugOperation(mod_5451_inner, "mod_5451");
    Operation_IFC mod_5452_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5452 <- mkDebugOperation(mod_5452_inner, "mod_5452");
    Operation_IFC mod_5453_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5453 <- mkDebugOperation(mod_5453_inner, "mod_5453");
    Operation_IFC mod_5454_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5454 <- mkDebugOperation(mod_5454_inner, "mod_5454");
    Operation_IFC mod_5455_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5455 <- mkDebugOperation(mod_5455_inner, "mod_5455");
    Operation_IFC mod_5456_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5456 <- mkDebugOperation(mod_5456_inner, "mod_5456");
    Operation_IFC mod_5457_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5457 <- mkDebugOperation(mod_5457_inner, "mod_5457");
    Operation_IFC mod_5458_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5458 <- mkDebugOperation(mod_5458_inner, "mod_5458");
    Operation_IFC mod_5459_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5459 <- mkDebugOperation(mod_5459_inner, "mod_5459");
    Operation_IFC mod_5460_inner <- mkRandomOffChipLoad(Cons(64, Cons(8, Cons(1, Cons(1, Cons(1, Cons(1, Nil)))))));
    Operation_IFC mod_5460 <- mkDebugOperation(mod_5460_inner, "mod_5460");
    Operation_IFC mod_5461_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5461 <- mkDebugOperation(mod_5461_inner, "mod_5461");
    Operation_IFC mod_5462_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5462 <- mkDebugOperation(mod_5462_inner, "mod_5462");
    Operation_IFC mod_5463_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5463 <- mkDebugOperation(mod_5463_inner, "mod_5463");
    Operation_IFC mod_5464_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5464 <- mkDebugOperation(mod_5464_inner, "mod_5464");
    Operation_IFC mod_5465_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5465 <- mkDebugOperation(mod_5465_inner, "mod_5465");
    Operation_IFC mod_5466_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5466 <- mkDebugOperation(mod_5466_inner, "mod_5466");
    Operation_IFC mod_5467_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5467 <- mkDebugOperation(mod_5467_inner, "mod_5467");
    Operation_IFC mod_5468_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5468 <- mkDebugOperation(mod_5468_inner, "mod_5468");
    Operation_IFC mod_5469_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5469 <- mkDebugOperation(mod_5469_inner, "mod_5469");
    Operation_IFC mod_5470_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5470 <- mkDebugOperation(mod_5470_inner, "mod_5470");
    Operation_IFC mod_5471_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5471 <- mkDebugOperation(mod_5471_inner, "mod_5471");
    Operation_IFC mod_5472_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5472 <- mkDebugOperation(mod_5472_inner, "mod_5472");
    Operation_IFC mod_5473_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5473 <- mkDebugOperation(mod_5473_inner, "mod_5473");
    Operation_IFC mod_5474_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5474 <- mkDebugOperation(mod_5474_inner, "mod_5474");
    Operation_IFC mod_5475_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5475 <- mkDebugOperation(mod_5475_inner, "mod_5475");
    Operation_IFC mod_5476_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5476 <- mkDebugOperation(mod_5476_inner, "mod_5476");
    Operation_IFC mod_5477_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5477 <- mkDebugOperation(mod_5477_inner, "mod_5477");
    Operation_IFC mod_5478_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5478 <- mkDebugOperation(mod_5478_inner, "mod_5478");
    Operation_IFC mod_5479_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5479 <- mkDebugOperation(mod_5479_inner, "mod_5479");
    Operation_IFC mod_5480_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5480 <- mkDebugOperation(mod_5480_inner, "mod_5480");
    Operation_IFC mod_5481_inner <- mkRandomSelectGen;
    Operation_IFC mod_5481 <- mkDebugOperation(mod_5481_inner, "mod_5481");
    Operation_IFC mod_5482_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5482 <- mkDebugOperation(mod_5482_inner, "mod_5482");
    Operation_IFC mod_5483_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5483 <- mkDebugOperation(mod_5483_inner, "mod_5483");
    Operation_IFC mod_5484_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5484 <- mkDebugOperation(mod_5484_inner, "mod_5484");
    Operation_IFC mod_5485_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5485 <- mkDebugOperation(mod_5485_inner, "mod_5485");
    Operation_IFC mod_5486_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5486 <- mkDebugOperation(mod_5486_inner, "mod_5486");
    Operation_IFC mod_5487_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5487 <- mkDebugOperation(mod_5487_inner, "mod_5487");
    Operation_IFC mod_5488_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5488 <- mkDebugOperation(mod_5488_inner, "mod_5488");
    Operation_IFC mod_5489_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5489 <- mkDebugOperation(mod_5489_inner, "mod_5489");
    Operation_IFC mod_5490_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5490 <- mkDebugOperation(mod_5490_inner, "mod_5490");
    Operation_IFC mod_5491_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5491 <- mkDebugOperation(mod_5491_inner, "mod_5491");
    Operation_IFC mod_5492_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5492 <- mkDebugOperation(mod_5492_inner, "mod_5492");
    Operation_IFC mod_5493_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5493 <- mkDebugOperation(mod_5493_inner, "mod_5493");
    Operation_IFC mod_5494_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5494 <- mkDebugOperation(mod_5494_inner, "mod_5494");
    Operation_IFC mod_5495_inner <- mkReshape(2, 1);
    Operation_IFC mod_5495 <- mkDebugOperation(mod_5495_inner, "mod_5495");
    Operation_IFC mod_5496_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5496 <- mkDebugOperation(mod_5496_inner, "mod_5496");
    Operation_IFC mod_5497_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5497 <- mkDebugOperation(mod_5497_inner, "mod_5497");
    Operation_IFC mod_5498_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5498 <- mkDebugOperation(mod_5498_inner, "mod_5498");
    Operation_IFC mod_5499_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5499 <- mkDebugOperation(mod_5499_inner, "mod_5499");
    Operation_IFC mod_5500_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5500 <- mkDebugOperation(mod_5500_inner, "mod_5500");
    Operation_IFC mod_5501_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5501 <- mkDebugOperation(mod_5501_inner, "mod_5501");
    Operation_IFC mod_5502_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5502 <- mkDebugOperation(mod_5502_inner, "mod_5502");
    Operation_IFC mod_5503_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5503 <- mkDebugOperation(mod_5503_inner, "mod_5503");
    Operation_IFC mod_5504_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5504 <- mkDebugOperation(mod_5504_inner, "mod_5504");
    Operation_IFC mod_5505_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5505 <- mkDebugOperation(mod_5505_inner, "mod_5505");
    Operation_IFC mod_5506_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5506 <- mkDebugOperation(mod_5506_inner, "mod_5506");
    Operation_IFC mod_5507_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5507 <- mkDebugOperation(mod_5507_inner, "mod_5507");
    Operation_IFC mod_5508_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5508 <- mkDebugOperation(mod_5508_inner, "mod_5508");
    Operation_IFC mod_5509_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5509 <- mkDebugOperation(mod_5509_inner, "mod_5509");
    Operation_IFC mod_5510_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5510 <- mkDebugOperation(mod_5510_inner, "mod_5510");
    Operation_IFC mod_5511_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5511 <- mkDebugOperation(mod_5511_inner, "mod_5511");
    Operation_IFC mod_5512_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5512 <- mkDebugOperation(mod_5512_inner, "mod_5512");
    Operation_IFC mod_5513_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5513 <- mkDebugOperation(mod_5513_inner, "mod_5513");
    Operation_IFC mod_5514_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5514 <- mkDebugOperation(mod_5514_inner, "mod_5514");
    Operation_IFC mod_5515_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5515 <- mkDebugOperation(mod_5515_inner, "mod_5515");
    Operation_IFC mod_5516_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5516 <- mkDebugOperation(mod_5516_inner, "mod_5516");
    Operation_IFC mod_5517_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5517 <- mkDebugOperation(mod_5517_inner, "mod_5517");
    Operation_IFC mod_5518_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5518 <- mkDebugOperation(mod_5518_inner, "mod_5518");
    Operation_IFC mod_5519_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5519 <- mkDebugOperation(mod_5519_inner, "mod_5519");
    Operation_IFC mod_5520_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5520 <- mkDebugOperation(mod_5520_inner, "mod_5520");
    Operation_IFC mod_5521_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5521 <- mkDebugOperation(mod_5521_inner, "mod_5521");
    Operation_IFC mod_5522_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5522 <- mkDebugOperation(mod_5522_inner, "mod_5522");
    Operation_IFC mod_5523_inner <- mkRepeatStatic(1);
    Operation_IFC mod_5523 <- mkDebugOperation(mod_5523_inner, "mod_5523");
    Operation_IFC mod_5524_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5524 <- mkDebugOperation(mod_5524_inner, "mod_5524");
    Operation_IFC mod_5525_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5525 <- mkDebugOperation(mod_5525_inner, "mod_5525");
    Operation_IFC mod_5526_inner <- mkRepeatStatic(1);
    Operation_IFC mod_5526 <- mkDebugOperation(mod_5526_inner, "mod_5526");
    Operation_IFC mod_5527_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5527 <- mkDebugOperation(mod_5527_inner, "mod_5527");
    Operation_IFC mod_5528_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5528 <- mkDebugOperation(mod_5528_inner, "mod_5528");
    Operation_IFC mod_5529_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5529 <- mkDebugOperation(mod_5529_inner, "mod_5529");
    Operation_IFC mod_5530_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5530 <- mkDebugOperation(mod_5530_inner, "mod_5530");
    Operation_IFC mod_5531_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5531 <- mkDebugOperation(mod_5531_inner, "mod_5531");
    Operation_IFC mod_5532_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5532 <- mkDebugOperation(mod_5532_inner, "mod_5532");
    Operation_IFC mod_5533_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5533 <- mkDebugOperation(mod_5533_inner, "mod_5533");
    Operation_IFC mod_5534_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5534 <- mkDebugOperation(mod_5534_inner, "mod_5534");
    Operation_IFC mod_5535_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5535 <- mkDebugOperation(mod_5535_inner, "mod_5535");
    Operation_IFC mod_5536_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5536 <- mkDebugOperation(mod_5536_inner, "mod_5536");
    Operation_IFC mod_5537_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5537 <- mkDebugOperation(mod_5537_inner, "mod_5537");
    Operation_IFC mod_5538_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5538 <- mkDebugOperation(mod_5538_inner, "mod_5538");
    Operation_IFC mod_5539_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5539 <- mkDebugOperation(mod_5539_inner, "mod_5539");
    Operation_IFC mod_5540_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5540 <- mkDebugOperation(mod_5540_inner, "mod_5540");
    Operation_IFC mod_5541_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5541 <- mkDebugOperation(mod_5541_inner, "mod_5541");
    Operation_IFC mod_5542_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5542 <- mkDebugOperation(mod_5542_inner, "mod_5542");
    Operation_IFC mod_5543_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5543 <- mkDebugOperation(mod_5543_inner, "mod_5543");
    Operation_IFC mod_5544_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5544 <- mkDebugOperation(mod_5544_inner, "mod_5544");
    Operation_IFC mod_5545_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5545 <- mkDebugOperation(mod_5545_inner, "mod_5545");
    Operation_IFC mod_5546_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5546 <- mkDebugOperation(mod_5546_inner, "mod_5546");
    Operation_IFC mod_5547_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5547 <- mkDebugOperation(mod_5547_inner, "mod_5547");
    Operation_IFC mod_5548_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5548 <- mkDebugOperation(mod_5548_inner, "mod_5548");
    Operation_IFC mod_5549_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5549 <- mkDebugOperation(mod_5549_inner, "mod_5549");
    Operation_IFC mod_5550_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5550 <- mkDebugOperation(mod_5550_inner, "mod_5550");
    Operation_IFC mod_5551_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5551 <- mkDebugOperation(mod_5551_inner, "mod_5551");
    Operation_IFC mod_5552_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5552 <- mkDebugOperation(mod_5552_inner, "mod_5552");
    Operation_IFC mod_5553_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5553 <- mkDebugOperation(mod_5553_inner, "mod_5553");
    Operation_IFC mod_5554_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5554 <- mkDebugOperation(mod_5554_inner, "mod_5554");
    Operation_IFC mod_5555_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5555 <- mkDebugOperation(mod_5555_inner, "mod_5555");
    Operation_IFC mod_5556_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5556 <- mkDebugOperation(mod_5556_inner, "mod_5556");
    Operation_IFC mod_5557_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5557 <- mkDebugOperation(mod_5557_inner, "mod_5557");
    Operation_IFC mod_5558_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5558 <- mkDebugOperation(mod_5558_inner, "mod_5558");
    Operation_IFC mod_5559_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5559 <- mkDebugOperation(mod_5559_inner, "mod_5559");
    Operation_IFC mod_5560_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5560 <- mkDebugOperation(mod_5560_inner, "mod_5560");
    Operation_IFC mod_5561_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5561 <- mkDebugOperation(mod_5561_inner, "mod_5561");
    Operation_IFC mod_5562_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5562 <- mkDebugOperation(mod_5562_inner, "mod_5562");
    Operation_IFC mod_5563_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5563 <- mkDebugOperation(mod_5563_inner, "mod_5563");
    Operation_IFC mod_5564_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5564 <- mkDebugOperation(mod_5564_inner, "mod_5564");
    Operation_IFC mod_5565_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5565 <- mkDebugOperation(mod_5565_inner, "mod_5565");
    Operation_IFC mod_5566_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5566 <- mkDebugOperation(mod_5566_inner, "mod_5566");
    Operation_IFC mod_5567_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5567 <- mkDebugOperation(mod_5567_inner, "mod_5567");
    Operation_IFC mod_5568_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5568 <- mkDebugOperation(mod_5568_inner, "mod_5568");
    Operation_IFC mod_5569_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5569 <- mkDebugOperation(mod_5569_inner, "mod_5569");
    Operation_IFC mod_5570_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5570 <- mkDebugOperation(mod_5570_inner, "mod_5570");
    Operation_IFC mod_5571_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5571 <- mkDebugOperation(mod_5571_inner, "mod_5571");
    Operation_IFC mod_5572_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5572 <- mkDebugOperation(mod_5572_inner, "mod_5572");
    Operation_IFC mod_5573_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5573 <- mkDebugOperation(mod_5573_inner, "mod_5573");
    Operation_IFC mod_5574_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5574 <- mkDebugOperation(mod_5574_inner, "mod_5574");
    Operation_IFC mod_5575_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5575 <- mkDebugOperation(mod_5575_inner, "mod_5575");
    Operation_IFC mod_5576_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5576 <- mkDebugOperation(mod_5576_inner, "mod_5576");
    Operation_IFC mod_5577_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5577 <- mkDebugOperation(mod_5577_inner, "mod_5577");
    Operation_IFC mod_5578_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5578 <- mkDebugOperation(mod_5578_inner, "mod_5578");
    Operation_IFC mod_5579_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5579 <- mkDebugOperation(mod_5579_inner, "mod_5579");
    Operation_IFC mod_5580_inner <- mkFlatten(1);
    Operation_IFC mod_5580 <- mkDebugOperation(mod_5580_inner, "mod_5580");
    Operation_IFC mod_5581_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5581 <- mkDebugOperation(mod_5581_inner, "mod_5581");
    Operation_IFC mod_5582_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5582 <- mkDebugOperation(mod_5582_inner, "mod_5582");
    Operation_IFC mod_5583_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5583 <- mkDebugOperation(mod_5583_inner, "mod_5583");
    Operation_IFC mod_5584_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5584 <- mkDebugOperation(mod_5584_inner, "mod_5584");
    Operation_IFC mod_5585_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5585 <- mkDebugOperation(mod_5585_inner, "mod_5585");
    Operation_IFC mod_5586_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5586 <- mkDebugOperation(mod_5586_inner, "mod_5586");
    Operation_IFC mod_5587_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5587 <- mkDebugOperation(mod_5587_inner, "mod_5587");
    Operation_IFC mod_5588_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5588 <- mkDebugOperation(mod_5588_inner, "mod_5588");
    Operation_IFC mod_5589_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5589 <- mkDebugOperation(mod_5589_inner, "mod_5589");
    Operation_IFC mod_5590_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5590 <- mkDebugOperation(mod_5590_inner, "mod_5590");
    Operation_IFC mod_5591_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5591 <- mkDebugOperation(mod_5591_inner, "mod_5591");
    Operation_IFC mod_5592_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5592 <- mkDebugOperation(mod_5592_inner, "mod_5592");
    Operation_IFC mod_5593_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5593 <- mkDebugOperation(mod_5593_inner, "mod_5593");
    Operation_IFC mod_5594_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5594 <- mkDebugOperation(mod_5594_inner, "mod_5594");
    Operation_IFC mod_5595_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5595 <- mkDebugOperation(mod_5595_inner, "mod_5595");
    Operation_IFC mod_5596_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5596 <- mkDebugOperation(mod_5596_inner, "mod_5596");
    Operation_IFC mod_5597_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5597 <- mkDebugOperation(mod_5597_inner, "mod_5597");
    Operation_IFC mod_5598_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5598 <- mkDebugOperation(mod_5598_inner, "mod_5598");
    Operation_IFC mod_5599_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5599 <- mkDebugOperation(mod_5599_inner, "mod_5599");
    Partition_IFC#(128) mod_5600_inner <- mkPartition(0, 128);
    Operation_IFC mod_5600 <- mkDebugOperation(mod_5600_inner.op, "mod_5600");
    Operation_IFC mod_5601_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5601 <- mkDebugOperation(mod_5601_inner, "mod_5601");
    Operation_IFC mod_5602_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5602 <- mkDebugOperation(mod_5602_inner, "mod_5602");
    Operation_IFC mod_5603_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5603 <- mkDebugOperation(mod_5603_inner, "mod_5603");
    Operation_IFC mod_5604_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5604 <- mkDebugOperation(mod_5604_inner, "mod_5604");
    Operation_IFC mod_5605_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5605 <- mkDebugOperation(mod_5605_inner, "mod_5605");
    Operation_IFC mod_5606_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5606 <- mkDebugOperation(mod_5606_inner, "mod_5606");
    Operation_IFC mod_5607_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5607 <- mkDebugOperation(mod_5607_inner, "mod_5607");
    Operation_IFC mod_5608_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5608 <- mkDebugOperation(mod_5608_inner, "mod_5608");
    Operation_IFC mod_5609_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5609 <- mkDebugOperation(mod_5609_inner, "mod_5609");
    Operation_IFC mod_5610_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5610 <- mkDebugOperation(mod_5610_inner, "mod_5610");
    Operation_IFC mod_5611_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5611 <- mkDebugOperation(mod_5611_inner, "mod_5611");
    Operation_IFC mod_5612_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5612 <- mkDebugOperation(mod_5612_inner, "mod_5612");
    Operation_IFC mod_5613_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5613 <- mkDebugOperation(mod_5613_inner, "mod_5613");
    Operation_IFC mod_5614_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5614 <- mkDebugOperation(mod_5614_inner, "mod_5614");
    Operation_IFC mod_5615_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5615 <- mkDebugOperation(mod_5615_inner, "mod_5615");
    Operation_IFC mod_5616_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5616 <- mkDebugOperation(mod_5616_inner, "mod_5616");
    Operation_IFC mod_5617_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5617 <- mkDebugOperation(mod_5617_inner, "mod_5617");
    Operation_IFC mod_5618_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5618 <- mkDebugOperation(mod_5618_inner, "mod_5618");
    Operation_IFC mod_5619_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5619 <- mkDebugOperation(mod_5619_inner, "mod_5619");
    Operation_IFC mod_5620_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5620 <- mkDebugOperation(mod_5620_inner, "mod_5620");
    Operation_IFC mod_5621_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5621 <- mkDebugOperation(mod_5621_inner, "mod_5621");
    Operation_IFC mod_5622_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5622 <- mkDebugOperation(mod_5622_inner, "mod_5622");
    Operation_IFC mod_5623_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5623 <- mkDebugOperation(mod_5623_inner, "mod_5623");
    Operation_IFC mod_5624_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5624 <- mkDebugOperation(mod_5624_inner, "mod_5624");
    Operation_IFC mod_5625_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5625 <- mkDebugOperation(mod_5625_inner, "mod_5625");
    Operation_IFC mod_5626_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5626 <- mkDebugOperation(mod_5626_inner, "mod_5626");
    Operation_IFC mod_5627_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5627 <- mkDebugOperation(mod_5627_inner, "mod_5627");
    Operation_IFC mod_5628_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5628 <- mkDebugOperation(mod_5628_inner, "mod_5628");
    Operation_IFC mod_5629_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5629 <- mkDebugOperation(mod_5629_inner, "mod_5629");
    Operation_IFC mod_5630_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5630 <- mkDebugOperation(mod_5630_inner, "mod_5630");
    Operation_IFC mod_5631_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5631 <- mkDebugOperation(mod_5631_inner, "mod_5631");
    Operation_IFC mod_5632_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5632 <- mkDebugOperation(mod_5632_inner, "mod_5632");
    Operation_IFC mod_5633_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5633 <- mkDebugOperation(mod_5633_inner, "mod_5633");
    Operation_IFC mod_5634_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5634 <- mkDebugOperation(mod_5634_inner, "mod_5634");
    Operation_IFC mod_5635_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5635 <- mkDebugOperation(mod_5635_inner, "mod_5635");
    Operation_IFC mod_5636_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5636 <- mkDebugOperation(mod_5636_inner, "mod_5636");
    Operation_IFC mod_5637_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5637 <- mkDebugOperation(mod_5637_inner, "mod_5637");
    Operation_IFC mod_5638_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5638 <- mkDebugOperation(mod_5638_inner, "mod_5638");
    Operation_IFC mod_5639_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5639 <- mkDebugOperation(mod_5639_inner, "mod_5639");
    Operation_IFC mod_5640_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5640 <- mkDebugOperation(mod_5640_inner, "mod_5640");
    Operation_IFC mod_5641_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5641 <- mkDebugOperation(mod_5641_inner, "mod_5641");
    Operation_IFC mod_5642_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5642 <- mkDebugOperation(mod_5642_inner, "mod_5642");
    Operation_IFC mod_5643_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5643 <- mkDebugOperation(mod_5643_inner, "mod_5643");
    Operation_IFC mod_5644_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5644 <- mkDebugOperation(mod_5644_inner, "mod_5644");
    Operation_IFC mod_5645_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5645 <- mkDebugOperation(mod_5645_inner, "mod_5645");
    Operation_IFC mod_5646_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5646 <- mkDebugOperation(mod_5646_inner, "mod_5646");
    Operation_IFC mod_5647_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5647 <- mkDebugOperation(mod_5647_inner, "mod_5647");
    Operation_IFC mod_5648_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5648 <- mkDebugOperation(mod_5648_inner, "mod_5648");
    (* descending_urgency = "rule_1, rule_2, rule_3, rule_4, rule_5, rule_6, rule_7, rule_8, rule_9, rule_10, rule_11, rule_12, rule_13, rule_14, rule_15, rule_16, rule_17, rule_18, rule_19, rule_20, rule_21, rule_22, rule_23, rule_24, rule_25, rule_26, rule_27, rule_28, rule_29, rule_30, rule_31, rule_32, rule_33, rule_34, rule_35, rule_36, rule_37, rule_38, rule_39, rule_40, rule_41, rule_42, rule_43, rule_44, rule_45, rule_46, rule_47, rule_48, rule_49, rule_50, rule_51, rule_52, rule_53, rule_54, rule_55, rule_56, rule_57, rule_58, rule_59, rule_60, rule_61, rule_62, rule_63, rule_64, rule_65, rule_66, rule_67, rule_68, rule_69, rule_70, rule_71, rule_72, rule_73, rule_74, rule_75, rule_76, rule_77, rule_78, rule_79, rule_80, rule_81, rule_82, rule_83, rule_84, rule_85, rule_86, rule_87, rule_88, rule_89, rule_90, rule_91, rule_92, rule_93, rule_94, rule_95, rule_96, rule_97, rule_98, rule_99, rule_100, rule_101, rule_102, rule_103, rule_104, rule_105, rule_106, rule_107, rule_108, rule_109, rule_110, rule_111, rule_112, rule_113, rule_114, rule_115, rule_116, rule_117, rule_118, rule_119, rule_120, rule_121, rule_122, rule_123, rule_124, rule_125, rule_126, rule_127, rule_128, rule_129, rule_130, rule_131, rule_132, rule_133, rule_134, rule_135, rule_136, rule_137, rule_138, rule_139, rule_140, rule_141, rule_142, rule_143, rule_144, rule_145, rule_146, rule_147, rule_148, rule_149, rule_150, rule_151, rule_152, rule_153, rule_154, rule_155, rule_156, rule_157, rule_158, rule_159, rule_160, rule_161, rule_162, rule_163, rule_164, rule_165, rule_166, rule_167, rule_168, rule_169, rule_170, rule_171, rule_172, rule_173, rule_174, rule_175, rule_176, rule_177, rule_178, rule_179, rule_180, rule_181, rule_182, rule_183, rule_184, rule_185, rule_186, rule_187, rule_188, rule_189, rule_190, rule_191, rule_192, rule_193, rule_194, rule_195, rule_196, rule_197, rule_198, rule_199, rule_200, rule_201, rule_202, rule_203, rule_204, rule_205, rule_206, rule_207, rule_208, rule_209, rule_210, rule_211, rule_212, rule_213, rule_214, rule_215, rule_216, rule_217, rule_218, rule_219, rule_220, rule_221, rule_222, rule_223, rule_224, rule_225, rule_226, rule_227, rule_228, rule_229, rule_230, rule_231, rule_232, rule_233, rule_234, rule_235, rule_236, rule_237, rule_238, rule_239, rule_240, rule_241, rule_242, rule_243, rule_244, rule_245, rule_246, rule_247, rule_248, rule_249, rule_250, rule_251, rule_252, rule_253, rule_254, rule_255, rule_256, rule_257, rule_258, rule_259, rule_260, rule_261, rule_262, rule_263, rule_264, rule_265, rule_266, rule_267, rule_268, rule_269, rule_270, rule_271, rule_272, rule_273, rule_274, rule_275, rule_276, rule_277, rule_278, rule_279, rule_280, rule_281, rule_282, rule_283, rule_284, rule_285, rule_286, rule_287, rule_288, rule_289, rule_290, rule_291, rule_292, rule_293, rule_294, rule_295, rule_296, rule_297, rule_298, rule_299, rule_300, rule_301, rule_302, rule_303, rule_304, rule_305, rule_306, rule_307, rule_308, rule_309, rule_310, rule_311, rule_312, rule_313, rule_314, rule_315, rule_316, rule_317, rule_318, rule_319, rule_320, rule_321, rule_322, rule_323, rule_324, rule_325, rule_326, rule_327, rule_328, rule_329, rule_330, rule_331, rule_332, rule_333, rule_334, rule_335, rule_336, rule_337, rule_338, rule_339, rule_340, rule_341, rule_342, rule_343, rule_344, rule_345, rule_346, rule_347, rule_348, rule_349, rule_350, rule_351, rule_352, rule_353, rule_354, rule_355, rule_356, rule_357, rule_358, rule_359, rule_360, rule_361, rule_362, rule_363, rule_364, rule_365, rule_366, rule_367, rule_368, rule_369, rule_370, rule_371, rule_372, rule_373, rule_374, rule_375, rule_376, rule_377, rule_378, rule_379, rule_380, rule_381, rule_382, rule_383, rule_384, rule_385, rule_386, rule_387, rule_388, rule_389, rule_390, rule_391, rule_392, rule_393, rule_394, rule_395, rule_396, rule_397, rule_398, rule_399, rule_400, rule_401, rule_402, rule_403, rule_404, rule_405, rule_406, rule_407, rule_408, rule_409, rule_410, rule_411, rule_412, rule_413, rule_414, rule_415, rule_416, rule_417, rule_418, rule_419, rule_420, rule_421, rule_422, rule_423, rule_424, rule_425, rule_426, rule_427, rule_428, rule_429, rule_430, rule_431, rule_432, rule_433, rule_434, rule_435, rule_436, rule_437, rule_438, rule_439, rule_440, rule_441, rule_442, rule_443, rule_444, rule_445, rule_446, rule_447, rule_448, rule_449, rule_450, rule_451, rule_452, rule_453, rule_454, rule_455, rule_456, rule_457, rule_458, rule_459, rule_460, rule_461, rule_462, rule_463, rule_464, rule_465, rule_466, rule_467, rule_468, rule_469, rule_470, rule_471, rule_472, rule_473, rule_474, rule_475, rule_476, rule_477, rule_478, rule_479, rule_480, rule_481, rule_482, rule_483, rule_484, rule_485, rule_486, rule_487, rule_488, rule_489, rule_490, rule_491, rule_492, rule_493, rule_494, rule_495, rule_496, rule_497, rule_498, rule_499, rule_500, rule_501, rule_502, rule_503, rule_504, rule_505, rule_506, rule_507, rule_508, rule_509, rule_510, rule_511, rule_512, rule_513, rule_514, rule_515, rule_516, rule_517, rule_518, rule_519, rule_520, rule_521, rule_522, rule_523, rule_524, rule_525, rule_526, rule_527, rule_528, rule_529, rule_530, rule_531, rule_532, rule_533, rule_534, rule_535, rule_536, rule_537, rule_538, rule_539, rule_540, rule_541, rule_542, rule_543, rule_544, rule_545, rule_546, rule_547, rule_548, rule_549, rule_550, rule_551, rule_552, rule_553, rule_554, rule_555, rule_556, rule_557, rule_558, rule_559, rule_560, rule_561, rule_562, rule_563, rule_564, rule_565, rule_566, rule_567, rule_568, rule_569, rule_570, rule_571, rule_572, rule_573, rule_574, rule_575, rule_576, rule_577, rule_578, rule_579, rule_580, rule_581, rule_582, rule_583, rule_584, rule_585, rule_586, rule_587, rule_588, rule_589, rule_590, rule_591, rule_592, rule_593, rule_594, rule_595, rule_596, rule_597, rule_598, rule_599, rule_600, rule_601, rule_602, rule_603, rule_604, rule_605, rule_606, rule_607, rule_608, rule_609, rule_610, rule_611, rule_612, rule_613, rule_614, rule_615, rule_616, rule_617, rule_618, rule_619, rule_620, rule_621, rule_622, rule_623, rule_624, rule_625, rule_626, rule_627, rule_628, rule_629, rule_630, rule_631, rule_632, rule_633, rule_634, rule_635, rule_636, rule_637, rule_638, rule_639, rule_640, rule_641, rule_642, rule_643, rule_644, rule_645, rule_646, rule_647, rule_648, rule_649, rule_650, rule_651, rule_652, rule_653, rule_654, rule_655, rule_656, rule_657, rule_658, rule_659, rule_660, rule_661, rule_662, rule_663, rule_664, rule_665, rule_666, rule_667, rule_668, rule_669, rule_670, rule_671, rule_672, rule_673, rule_674, rule_675, rule_676, rule_677, rule_678, rule_679, rule_680, rule_681, rule_682, rule_683, rule_684, rule_685, rule_686, rule_687, rule_688, rule_689, rule_690, rule_691, rule_692, rule_693, rule_694, rule_695, rule_696, rule_697, rule_698, rule_699, rule_700, rule_701, rule_702, rule_703, rule_704, rule_705, rule_706, rule_707, rule_708, rule_709, rule_710, rule_711, rule_712, rule_713, rule_714, rule_715, rule_716, rule_717, rule_718, rule_719, rule_720, rule_721, rule_722, rule_723, rule_724, rule_725, rule_726, rule_727, rule_728, rule_729, rule_730, rule_731, rule_732, rule_733, rule_734, rule_735, rule_736, rule_737, rule_738, rule_739, rule_740, rule_741, rule_742, rule_743, rule_744, rule_745, rule_746, rule_747, rule_748, rule_749, rule_750, rule_751, rule_752, rule_753, rule_754, rule_755, rule_756, rule_757, rule_758, rule_759, rule_760, rule_761, rule_762, rule_763, rule_764, rule_765, rule_766, rule_767, rule_768, rule_769, rule_770, rule_771, rule_772, rule_773, rule_774, rule_775, rule_776, rule_777, rule_778, rule_779, rule_780, rule_781, rule_782, rule_783, rule_784, rule_785, rule_786, rule_787, rule_788, rule_789, rule_790, rule_791, rule_792, rule_793, rule_794, rule_795, rule_796, rule_797, rule_798, rule_799, rule_800, rule_801, rule_802, rule_803, rule_804, rule_805, rule_806, rule_807, rule_808, rule_809, rule_810, rule_811, rule_812, rule_813, rule_814, rule_815, rule_816, rule_817, rule_818, rule_819, rule_820, rule_821, rule_822, rule_823, rule_824, rule_825, rule_826, rule_827, rule_828, rule_829, rule_830, rule_831, rule_832, rule_833, rule_834, rule_835, rule_836, rule_837, rule_838, rule_839, rule_840, rule_841, rule_842, rule_843, rule_844, rule_845, rule_846, rule_847, rule_848, rule_849, rule_850, rule_851, rule_852, rule_853, rule_854, rule_855, rule_856, rule_857, rule_858, rule_859, rule_860, rule_861, rule_862, rule_863, rule_864, rule_865, rule_866, rule_867, rule_868, rule_869, rule_870, rule_871, rule_872, rule_873, rule_874, rule_875, rule_876, rule_877, rule_878, rule_879, rule_880, rule_881, rule_882, rule_883, rule_884, rule_885, rule_886, rule_887, rule_888, rule_889, rule_890, rule_891, rule_892, rule_893, rule_894, rule_895, rule_896, rule_897, rule_898, rule_899, rule_900, rule_901, rule_902, rule_903, rule_904, rule_905, rule_906, rule_907, rule_908, rule_909, rule_910, rule_911, rule_912, rule_913, rule_914, rule_915, rule_916, rule_917, rule_918, rule_919, rule_920, rule_921, rule_922, rule_923, rule_924, rule_925, rule_926, rule_927, rule_928, rule_929, rule_930, rule_931, rule_932, rule_933, rule_934, rule_935, rule_936, rule_937, rule_938, rule_939, rule_940, rule_941, rule_942, rule_943, rule_944, rule_945, rule_946, rule_947, rule_948, rule_949, rule_950, rule_951, rule_952, rule_953, rule_954, rule_955, rule_956, rule_957, rule_958, rule_959, rule_960, rule_961, rule_962, rule_963, rule_964, rule_965, rule_966, rule_967, rule_968, rule_969, rule_970, rule_971, rule_972, rule_973, rule_974, rule_975, rule_976, rule_977, rule_978, rule_979, rule_980, rule_981, rule_982, rule_983, rule_984, rule_985, rule_986, rule_987, rule_988, rule_989, rule_990, rule_991, rule_992, rule_993, rule_994, rule_995, rule_996, rule_997, rule_998, rule_999, rule_1000, rule_1001, rule_1002, rule_1003, rule_1004, rule_1005, rule_1006, rule_1007, rule_1008, rule_1009, rule_1010, rule_1011, rule_1012, rule_1013, rule_1014, rule_1015, rule_1016, rule_1017, rule_1018, rule_1019, rule_1020, rule_1021, rule_1022, rule_1023, rule_1024, rule_1025, rule_1026, rule_1027, rule_1028, rule_1029, rule_1030, rule_1031, rule_1032, rule_1033, rule_1034, rule_1035, rule_1036, rule_1037, rule_1038, rule_1039, rule_1040, rule_1041, rule_1042, rule_1043, rule_1044, rule_1045, rule_1046, rule_1047, rule_1048, rule_1049, rule_1050, rule_1051, rule_1052, rule_1053, rule_1054, rule_1055, rule_1056, rule_1057, rule_1058, rule_1059, rule_1060, rule_1061, rule_1062, rule_1063, rule_1064, rule_1065, rule_1066, rule_1067, rule_1068, rule_1069, rule_1070, rule_1071, rule_1072, rule_1073, rule_1074, rule_1075, rule_1076, rule_1077, rule_1078, rule_1079, rule_1080, rule_1081, rule_1082, rule_1083, rule_1084, rule_1085, rule_1086, rule_1087, rule_1088, rule_1089, rule_1090, rule_1091, rule_1092, rule_1093, rule_1094, rule_1095, rule_1096, rule_1097, rule_1098, rule_1099, rule_1100, rule_1101, rule_1102, rule_1103, rule_1104, rule_1105, rule_1106, rule_1107, rule_1108, rule_1109, rule_1110, rule_1111, rule_1112, rule_1113, rule_1114, rule_1115, rule_1116, rule_1117, rule_1118, rule_1119, rule_1120, rule_1121, rule_1122, rule_1123, rule_1124, rule_1125, rule_1126, rule_1127, rule_1128, rule_1129, rule_1130, rule_1131, rule_1132, rule_1133, rule_1134, rule_1135, rule_1136, rule_1137, rule_1138, rule_1139, rule_1140, rule_1141, rule_1142, rule_1143, rule_1144, rule_1145, rule_1146, rule_1147, rule_1148, rule_1149, rule_1150, rule_1151, rule_1152, rule_1153, rule_1154, rule_1155, rule_1156, rule_1157, rule_1158, rule_1159, rule_1160, rule_1161, rule_1162, rule_1163, rule_1164, rule_1165, rule_1166, rule_1167, rule_1168, rule_1169, rule_1170, rule_1171, rule_1172, rule_1173, rule_1174, rule_1175, rule_1176, rule_1177, rule_1178, rule_1179, rule_1180, rule_1181, rule_1182, rule_1183, rule_1184, rule_1185, rule_1186, rule_1187, rule_1188, rule_1189, rule_1190, rule_1191, rule_1192, rule_1193, rule_1194, rule_1195, rule_1196, rule_1197, rule_1198, rule_1199, rule_1200, rule_1201, rule_1202, rule_1203, rule_1204, rule_1205, rule_1206, rule_1207, rule_1208, rule_1209, rule_1210, rule_1211, rule_1212, rule_1213, rule_1214, rule_1215, rule_1216, rule_1217, rule_1218, rule_1219, rule_1220, rule_1221, rule_1222, rule_1223, rule_1224, rule_1225, rule_1226, rule_1227, rule_1228, rule_1229, rule_1230, rule_1231, rule_1232, rule_1233, rule_1234, rule_1235, rule_1236, rule_1237, rule_1238, rule_1239, rule_1240, rule_1241, rule_1242, rule_1243, rule_1244, rule_1245, rule_1246, rule_1247, rule_1248, rule_1249, rule_1250, rule_1251, rule_1252, rule_1253, rule_1254, rule_1255, rule_1256, rule_1257, rule_1258, rule_1259, rule_1260, rule_1261, rule_1262, rule_1263, rule_1264, rule_1265, rule_1266, rule_1267, rule_1268, rule_1269, rule_1270, rule_1271, rule_1272, rule_1273, rule_1274, rule_1275, rule_1276, rule_1277, rule_1278, rule_1279, rule_1280, rule_1281, rule_1282, rule_1283, rule_1284, rule_1285, rule_1286, rule_1287, rule_1288, rule_1289, rule_1290, rule_1291, rule_1292, rule_1293, rule_1294, rule_1295, rule_1296, rule_1297, rule_1298, rule_1299, rule_1300, rule_1301, rule_1302, rule_1303, rule_1304, rule_1305, rule_1306, rule_1307, rule_1308, rule_1309, rule_1310, rule_1311, rule_1312, rule_1313, rule_1314, rule_1315, rule_1316, rule_1317, rule_1318, rule_1319, rule_1320, rule_1321, rule_1322, rule_1323, rule_1324, rule_1325, rule_1326, rule_1327, rule_1328, rule_1329, rule_1330, rule_1331, rule_1332, rule_1333, rule_1334, rule_1335, rule_1336, rule_1337, rule_1338, rule_1339, rule_1340, rule_1341, rule_1342, rule_1343, rule_1344, rule_1345, rule_1346, rule_1347, rule_1348, rule_1349, rule_1350, rule_1351, rule_1352, rule_1353, rule_1354, rule_1355, rule_1356, rule_1357, rule_1358, rule_1359, rule_1360, rule_1361, rule_1362, rule_1363, rule_1364, rule_1365, rule_1366, rule_1367, rule_1368, rule_1369, rule_1370, rule_1371, rule_1372, rule_1373, rule_1374, rule_1375, rule_1376, rule_1377, rule_1378, rule_1379, rule_1380, rule_1381, rule_1382, rule_1383, rule_1384, rule_1385, rule_1386, rule_1387, rule_1388, rule_1389, rule_1390, rule_1391, rule_1392, rule_1393, rule_1394, rule_1395, rule_1396, rule_1397, rule_1398, rule_1399, rule_1400, rule_1401, rule_1402, rule_1403, rule_1404, rule_1405, rule_1406, rule_1407, rule_1408, rule_1409, rule_1410, rule_1411, rule_1412, rule_1413, rule_1414, rule_1415, rule_1416, rule_1417, rule_1418, rule_1419, rule_1420, rule_1421, rule_1422, rule_1423, rule_1424, rule_1425, rule_1426, rule_1427, rule_1428, rule_1429, rule_1430, rule_1431, rule_1432, rule_1433, rule_1434, rule_1435, rule_1436, rule_1437, rule_1438, rule_1439, rule_1440, rule_1441, rule_1442, rule_1443, rule_1444, rule_1445, rule_1446, rule_1447, rule_1448, rule_1449, rule_1450, rule_1451, rule_1452, rule_1453, rule_1454, rule_1455, rule_1456, rule_1457, rule_1458, rule_1459, rule_1460, rule_1461, rule_1462, rule_1463, rule_1464, rule_1465, rule_1466, rule_1467, rule_1468, rule_1469, rule_1470, rule_1471, rule_1472, rule_1473, rule_1474, rule_1475, rule_1476, rule_1477, rule_1478, rule_1479, rule_1480, rule_1481, rule_1482, rule_1483, rule_1484, rule_1485, rule_1486, rule_1487, rule_1488, rule_1489, rule_1490, rule_1491, rule_1492, rule_1493, rule_1494, rule_1495, rule_1496, rule_1497, rule_1498, rule_1499, rule_1500, rule_1501, rule_1502, rule_1503, rule_1504, rule_1505, rule_1506, rule_1507, rule_1508, rule_1509, rule_1510, rule_1511, rule_1512, rule_1513, rule_1514, rule_1515, rule_1516, rule_1517, rule_1518, rule_1519, rule_1520, rule_1521, rule_1522, rule_1523, rule_1524, rule_1525, rule_1526, rule_1527, rule_1528, rule_1529, rule_1530, rule_1531, rule_1532, rule_1533, rule_1534, rule_1535, rule_1536, rule_1537, rule_1538, rule_1539, rule_1540, rule_1541, rule_1542, rule_1543, rule_1544, rule_1545, rule_1546, rule_1547, rule_1548, rule_1549, rule_1550, rule_1551, rule_1552, rule_1553, rule_1554, rule_1555, rule_1556, rule_1557, rule_1558, rule_1559, rule_1560, rule_1561, rule_1562, rule_1563, rule_1564, rule_1565, rule_1566, rule_1567, rule_1568, rule_1569, rule_1570, rule_1571, rule_1572, rule_1573, rule_1574, rule_1575, rule_1576, rule_1577, rule_1578, rule_1579, rule_1580, rule_1581, rule_1582, rule_1583, rule_1584, rule_1585, rule_1586, rule_1587, rule_1588, rule_1589, rule_1590, rule_1591, rule_1592, rule_1593, rule_1594, rule_1595, rule_1596, rule_1597, rule_1598, rule_1599, rule_1600, rule_1601, rule_1602, rule_1603, rule_1604, rule_1605, rule_1606, rule_1607, rule_1608, rule_1609, rule_1610, rule_1611, rule_1612, rule_1613, rule_1614, rule_1615, rule_1616, rule_1617, rule_1618, rule_1619, rule_1620, rule_1621, rule_1622, rule_1623, rule_1624, rule_1625, rule_1626, rule_1627, rule_1628, rule_1629, rule_1630, rule_1631, rule_1632, rule_1633, rule_1634, rule_1635, rule_1636, rule_1637, rule_1638, rule_1639, rule_1640, rule_1641, rule_1642, rule_1643, rule_1644, rule_1645, rule_1646, rule_1647, rule_1648, rule_1649, rule_1650, rule_1651, rule_1652, rule_1653, rule_1654, rule_1655, rule_1656, rule_1657, rule_1658, rule_1659, rule_1660, rule_1661, rule_1662, rule_1663, rule_1664, rule_1665, rule_1666, rule_1667, rule_1668, rule_1669, rule_1670, rule_1671, rule_1672, rule_1673, rule_1674, rule_1675, rule_1676, rule_1677, rule_1678, rule_1679, rule_1680, rule_1681, rule_1682, rule_1683, rule_1684, rule_1685, rule_1686, rule_1687, rule_1688, rule_1689, rule_1690, rule_1691, rule_1692, rule_1693, rule_1694, rule_1695, rule_1696, rule_1697, rule_1698, rule_1699, rule_1700, rule_1701, rule_1702, rule_1703, rule_1704, rule_1705, rule_1706, rule_1707, rule_1708, rule_1709, rule_1710, rule_1711, rule_1712, rule_1713, rule_1714, rule_1715, rule_1716, rule_1717, rule_1718, rule_1719, rule_1720, rule_1721, rule_1722, rule_1723, rule_1724, rule_1725, rule_1726, rule_1727, rule_1728, rule_1729, rule_1730, rule_1731, rule_1732, rule_1733, rule_1734, rule_1735, rule_1736, rule_1737, rule_1738, rule_1739, rule_1740, rule_1741, rule_1742, rule_1743, rule_1744, rule_1745, rule_1746, rule_1747, rule_1748, rule_1749, rule_1750, rule_1751, rule_1752, rule_1753, rule_1754, rule_1755, rule_1756, rule_1757, rule_1758, rule_1759, rule_1760, rule_1761, rule_1762, rule_1763, rule_1764, rule_1765, rule_1766, rule_1767, rule_1768, rule_1769, rule_1770, rule_1771, rule_1772, rule_1773, rule_1774, rule_1775, rule_1776, rule_1777, rule_1778, rule_1779, rule_1780, rule_1781, rule_1782, rule_1783, rule_1784, rule_1785, rule_1786, rule_1787, rule_1788, rule_1789, rule_1790, rule_1791, rule_1792, rule_1793, rule_1794, rule_1795, rule_1796, rule_1797, rule_1798, rule_1799, rule_1800, rule_1801, rule_1802, rule_1803, rule_1804, rule_1805, rule_1806, rule_1807, rule_1808, rule_1809, rule_1810, rule_1811, rule_1812, rule_1813, rule_1814, rule_1815, rule_1816, rule_1817, rule_1818, rule_1819, rule_1820, rule_1821, rule_1822, rule_1823, rule_1824, rule_1825, rule_1826, rule_1827, rule_1828, rule_1829, rule_1830, rule_1831, rule_1832, rule_1833, rule_1834, rule_1835, rule_1836, rule_1837, rule_1838, rule_1839, rule_1840, rule_1841, rule_1842, rule_1843, rule_1844, rule_1845, rule_1846, rule_1847, rule_1848, rule_1849, rule_1850, rule_1851, rule_1852, rule_1853, rule_1854, rule_1855, rule_1856, rule_1857, rule_1858, rule_1859, rule_1860, rule_1861, rule_1862, rule_1863, rule_1864, rule_1865, rule_1866, rule_1867, rule_1868, rule_1869, rule_1870, rule_1871, rule_1872, rule_1873, rule_1874, rule_1875, rule_1876, rule_1877, rule_1878, rule_1879, rule_1880, rule_1881, rule_1882, rule_1883, rule_1884, rule_1885, rule_1886, rule_1887, rule_1888, rule_1889, rule_1890, rule_1891, rule_1892, rule_1893, rule_1894, rule_1895, rule_1896, rule_1897, rule_1898, rule_1899, rule_1900, rule_1901, rule_1902, rule_1903, rule_1904, rule_1905, rule_1906, rule_1907, rule_1908, rule_1909, rule_1910, rule_1911, rule_1912, rule_1913, rule_1914, rule_1915, rule_1916, rule_1917, rule_1918, rule_1919, rule_1920, rule_1921, rule_1922, rule_1923, rule_1924, rule_1925, rule_1926, rule_1927, rule_1928, rule_1929, rule_1930, rule_1931, rule_1932, rule_1933, rule_1934, rule_1935, rule_1936, rule_1937, rule_1938, rule_1939, rule_1940, rule_1941, rule_1942, rule_1943, rule_1944, rule_1945, rule_1946, rule_1947, rule_1948, rule_1949, rule_1950, rule_1951, rule_1952, rule_1953, rule_1954, rule_1955, rule_1956, rule_1957, rule_1958, rule_1959, rule_1960, rule_1961, rule_1962, rule_1963, rule_1964, rule_1965, rule_1966, rule_1967, rule_1968, rule_1969, rule_1970, rule_1971, rule_1972, rule_1973, rule_1974, rule_1975, rule_1976, rule_1977, rule_1978, rule_1979, rule_1980, rule_1981, rule_1982, rule_1983, rule_1984, rule_1985, rule_1986, rule_1987, rule_1988, rule_1989, rule_1990, rule_1991, rule_1992, rule_1993, rule_1994, rule_1995, rule_1996, rule_1997, rule_1998, rule_1999, rule_2000, rule_2001, rule_2002, rule_2003, rule_2004, rule_2005, rule_2006, rule_2007, rule_2008, rule_2009, rule_2010, rule_2011, rule_2012, rule_2013, rule_2014, rule_2015, rule_2016, rule_2017, rule_2018, rule_2019, rule_2020, rule_2021, rule_2022, rule_2023, rule_2024, rule_2025, rule_2026, rule_2027, rule_2028, rule_2029, rule_2030, rule_2031, rule_2032, rule_2033, rule_2034, rule_2035, rule_2036, rule_2037, rule_2038, rule_2039, rule_2040, rule_2041, rule_2042, rule_2043, rule_2044, rule_2045, rule_2046, rule_2047, rule_2048, rule_2049, rule_2050, rule_2051, rule_2052, rule_2053, rule_2054, rule_2055, rule_2056, rule_2057, rule_2058, rule_2059, rule_2060, rule_2061, rule_2062, rule_2063, rule_2064, rule_2065, rule_2066, rule_2067, rule_2068, rule_2069, rule_2070, rule_2071, rule_2072, rule_2073, rule_2074, rule_2075, rule_2076, rule_2077, rule_2078, rule_2079, rule_2080, rule_2081, rule_2082, rule_2083, rule_2084, rule_2085, rule_2086, rule_2087, rule_2088, rule_2089, rule_2090, rule_2091, rule_2092, rule_2093, rule_2094, rule_2095, rule_2096, rule_2097, rule_2098, rule_2099, rule_2100, rule_2101, rule_2102, rule_2103, rule_2104, rule_2105, rule_2106, rule_2107, rule_2108, rule_2109, rule_2110, rule_2111, rule_2112, rule_2113, rule_2114, rule_2115, rule_2116, rule_2117, rule_2118, rule_2119, rule_2120, rule_2121, rule_2122, rule_2123, rule_2124, rule_2125, rule_2126, rule_2127, rule_2128, rule_2129, rule_2130, rule_2131, rule_2132, rule_2133, rule_2134, rule_2135, rule_2136, rule_2137, rule_2138, rule_2139, rule_2140, rule_2141, rule_2142, rule_2143, rule_2144, rule_2145, rule_2146, rule_2147, rule_2148, rule_2149, rule_2150, rule_2151, rule_2152, rule_2153, rule_2154, rule_2155, rule_2156, rule_2157, rule_2158, rule_2159, rule_2160, rule_2161, rule_2162, rule_2163, rule_2164, rule_2165, rule_2166, rule_2167, rule_2168, rule_2169, rule_2170, rule_2171, rule_2172, rule_2173, rule_2174, rule_2175, rule_2176, rule_2177, rule_2178, rule_2179, rule_2180, rule_2181, rule_2182, rule_2183, rule_2184, rule_2185, rule_2186, rule_2187, rule_2188, rule_2189, rule_2190, rule_2191, rule_2192, rule_2193, rule_2194, rule_2195, rule_2196, rule_2197, rule_2198, rule_2199, rule_2200, rule_2201, rule_2202, rule_2203, rule_2204, rule_2205, rule_2206, rule_2207, rule_2208, rule_2209, rule_2210, rule_2211, rule_2212, rule_2213, rule_2214, rule_2215, rule_2216, rule_2217, rule_2218, rule_2219, rule_2220, rule_2221, rule_2222, rule_2223, rule_2224, rule_2225, rule_2226, rule_2227, rule_2228, rule_2229, rule_2230, rule_2231, rule_2232, rule_2233, rule_2234, rule_2235, rule_2236, rule_2237, rule_2238, rule_2239, rule_2240, rule_2241, rule_2242, rule_2243, rule_2244, rule_2245, rule_2246, rule_2247, rule_2248, rule_2249, rule_2250, rule_2251, rule_2252, rule_2253, rule_2254, rule_2255, rule_2256, rule_2257, rule_2258, rule_2259, rule_2260, rule_2261, rule_2262, rule_2263, rule_2264, rule_2265, rule_2266, rule_2267, rule_2268, rule_2269, rule_2270, rule_2271, rule_2272, rule_2273, rule_2274, rule_2275, rule_2276, rule_2277, rule_2278, rule_2279, rule_2280, rule_2281, rule_2282, rule_2283, rule_2284, rule_2285, rule_2286, rule_2287, rule_2288, rule_2289, rule_2290, rule_2291, rule_2292, rule_2293, rule_2294, rule_2295, rule_2296, rule_2297, rule_2298, rule_2299, rule_2300, rule_2301, rule_2302, rule_2303, rule_2304, rule_2305, rule_2306, rule_2307, rule_2308, rule_2309, rule_2310, rule_2311, rule_2312, rule_2313, rule_2314, rule_2315, rule_2316, rule_2317, rule_2318, rule_2319, rule_2320, rule_2321, rule_2322, rule_2323, rule_2324, rule_2325, rule_2326, rule_2327, rule_2328, rule_2329, rule_2330, rule_2331, rule_2332, rule_2333, rule_2334, rule_2335, rule_2336, rule_2337, rule_2338, rule_2339, rule_2340, rule_2341, rule_2342, rule_2343, rule_2344, rule_2345, rule_2346, rule_2347, rule_2348, rule_2349, rule_2350, rule_2351, rule_2352, rule_2353, rule_2354, rule_2355, rule_2356, rule_2357, rule_2358, rule_2359, rule_2360, rule_2361, rule_2362, rule_2363, rule_2364, rule_2365, rule_2366, rule_2367, rule_2368, rule_2369, rule_2370, rule_2371, rule_2372, rule_2373, rule_2374, rule_2375, rule_2376, rule_2377, rule_2378, rule_2379, rule_2380, rule_2381, rule_2382, rule_2383, rule_2384, rule_2385, rule_2386, rule_2387, rule_2388, rule_2389, rule_2390, rule_2391, rule_2392, rule_2393, rule_2394, rule_2395, rule_2396, rule_2397, rule_2398, rule_2399, rule_2400, rule_2401, rule_2402, rule_2403, rule_2404, rule_2405, rule_2406, rule_2407, rule_2408, rule_2409, rule_2410, rule_2411, rule_2412, rule_2413, rule_2414, rule_2415, rule_2416, rule_2417, rule_2418, rule_2419, rule_2420, rule_2421, rule_2422, rule_2423, rule_2424, rule_2425, rule_2426, rule_2427, rule_2428, rule_2429, rule_2430, rule_2431, rule_2432, rule_2433, rule_2434, rule_2435, rule_2436, rule_2437, rule_2438, rule_2439, rule_2440, rule_2441, rule_2442, rule_2443, rule_2444, rule_2445, rule_2446, rule_2447, rule_2448, rule_2449, rule_2450, rule_2451, rule_2452, rule_2453, rule_2454, rule_2455, rule_2456, rule_2457, rule_2458, rule_2459, rule_2460, rule_2461, rule_2462, rule_2463, rule_2464, rule_2465, rule_2466, rule_2467, rule_2468, rule_2469, rule_2470, rule_2471, rule_2472, rule_2473, rule_2474, rule_2475, rule_2476, rule_2477, rule_2478, rule_2479, rule_2480, rule_2481, rule_2482, rule_2483, rule_2484, rule_2485, rule_2486, rule_2487, rule_2488, rule_2489, rule_2490, rule_2491, rule_2492, rule_2493, rule_2494, rule_2495, rule_2496, rule_2497, rule_2498, rule_2499, rule_2500, rule_2501, rule_2502, rule_2503, rule_2504, rule_2505, rule_2506, rule_2507, rule_2508, rule_2509, rule_2510, rule_2511, rule_2512, rule_2513, rule_2514, rule_2515, rule_2516, rule_2517, rule_2518, rule_2519, rule_2520, rule_2521, rule_2522, rule_2523, rule_2524, rule_2525, rule_2526, rule_2527, rule_2528, rule_2529, rule_2530, rule_2531, rule_2532, rule_2533, rule_2534, rule_2535, rule_2536, rule_2537, rule_2538, rule_2539, rule_2540, rule_2541, rule_2542, rule_2543, rule_2544, rule_2545, rule_2546, rule_2547, rule_2548, rule_2549, rule_2550, rule_2551, rule_2552, rule_2553, rule_2554, rule_2555, rule_2556, rule_2557, rule_2558, rule_2559, rule_2560, rule_2561, rule_2562, rule_2563, rule_2564, rule_2565, rule_2566, rule_2567, rule_2568, rule_2569, rule_2570, rule_2571, rule_2572, rule_2573, rule_2574, rule_2575, rule_2576, rule_2577, rule_2578, rule_2579, rule_2580, rule_2581, rule_2582, rule_2583, rule_2584, rule_2585, rule_2586, rule_2587, rule_2588, rule_2589, rule_2590, rule_2591, rule_2592, rule_2593, rule_2594, rule_2595, rule_2596, rule_2597, rule_2598, rule_2599, rule_2600, rule_2601, rule_2602, rule_2603, rule_2604, rule_2605, rule_2606, rule_2607, rule_2608, rule_2609, rule_2610, rule_2611, rule_2612, rule_2613, rule_2614, rule_2615, rule_2616, rule_2617, rule_2618, rule_2619, rule_2620, rule_2621, rule_2622, rule_2623, rule_2624, rule_2625, rule_2626, rule_2627, rule_2628, rule_2629, rule_2630, rule_2631, rule_2632, rule_2633, rule_2634, rule_2635, rule_2636, rule_2637, rule_2638, rule_2639, rule_2640, rule_2641, rule_2642, rule_2643, rule_2644, rule_2645, rule_2646, rule_2647, rule_2648, rule_2649, rule_2650, rule_2651, rule_2652, rule_2653, rule_2654, rule_2655, rule_2656, rule_2657, rule_2658, rule_2659, rule_2660, rule_2661, rule_2662, rule_2663, rule_2664, rule_2665, rule_2666, rule_2667, rule_2668, rule_2669, rule_2670, rule_2671, rule_2672, rule_2673, rule_2674, rule_2675, rule_2676, rule_2677, rule_2678, rule_2679, rule_2680, rule_2681, rule_2682, rule_2683, rule_2684, rule_2685, rule_2686, rule_2687, rule_2688, rule_2689, rule_2690, rule_2691, rule_2692, rule_2693, rule_2694, rule_2695, rule_2696, rule_2697, rule_2698, rule_2699, rule_2700, rule_2701, rule_2702, rule_2703, rule_2704, rule_2705, rule_2706, rule_2707, rule_2708, rule_2709, rule_2710, rule_2711, rule_2712, rule_2713, rule_2714, rule_2715, rule_2716, rule_2717, rule_2718, rule_2719, rule_2720, rule_2721, rule_2722, rule_2723, rule_2724, rule_2725, rule_2726, rule_2727, rule_2728, rule_2729, rule_2730, rule_2731, rule_2732, rule_2733, rule_2734, rule_2735, rule_2736, rule_2737, rule_2738, rule_2739, rule_2740, rule_2741, rule_2742, rule_2743, rule_2744, rule_2745, rule_2746, rule_2747, rule_2748, rule_2749, rule_2750, rule_2751, rule_2752, rule_2753, rule_2754, rule_2755, rule_2756, rule_2757, rule_2758, rule_2759, rule_2760, rule_2761, rule_2762, rule_2763, rule_2764, rule_2765, rule_2766, rule_2767, rule_2768, rule_2769, rule_2770, rule_2771, rule_2772, rule_2773, rule_2774, rule_2775, rule_2776, rule_2777, rule_2778, rule_2779, rule_2780, rule_2781, rule_2782, rule_2783, rule_2784, rule_2785, rule_2786, rule_2787, rule_2788, rule_2789, rule_2790, rule_2791, rule_2792, rule_2793, rule_2794, rule_2795, rule_2796, rule_2797, rule_2798, rule_2799, rule_2800, rule_2801, rule_2802, rule_2803, rule_2804, rule_2805, rule_2806, rule_2807, rule_2808, rule_2809, rule_2810, rule_2811, rule_2812, rule_2813, rule_2814, rule_2815, rule_2816, rule_2817, rule_2818, rule_2819, rule_2820, rule_2821, rule_2822, rule_2823, rule_2824, rule_2825, rule_2826, rule_2827, rule_2828, rule_2829, rule_2830, rule_2831, rule_2832, rule_2833, rule_2834, rule_2835, rule_2836, rule_2837, rule_2838, rule_2839, rule_2840, rule_2841, rule_2842, rule_2843, rule_2844, rule_2845, rule_2846, rule_2847, rule_2848, rule_2849, rule_2850, rule_2851, rule_2852, rule_2853, rule_2854, rule_2855, rule_2856, rule_2857, rule_2858, rule_2859, rule_2860, rule_2861, rule_2862, rule_2863, rule_2864, rule_2865, rule_2866, rule_2867, rule_2868, rule_2869, rule_2870, rule_2871, rule_2872, rule_2873, rule_2874, rule_2875, rule_2876, rule_2877, rule_2878, rule_2879, rule_2880, rule_2881, rule_2882, rule_2883, rule_2884, rule_2885, rule_2886, rule_2887, rule_2888, rule_2889, rule_2890, rule_2891, rule_2892, rule_2893, rule_2894, rule_2895, rule_2896, rule_2897, rule_2898, rule_2899, rule_2900, rule_2901, rule_2902, rule_2903, rule_2904, rule_2905, rule_2906, rule_2907, rule_2908, rule_2909, rule_2910, rule_2911, rule_2912, rule_2913, rule_2914, rule_2915, rule_2916, rule_2917, rule_2918, rule_2919, rule_2920, rule_2921, rule_2922, rule_2923, rule_2924, rule_2925, rule_2926, rule_2927, rule_2928, rule_2929, rule_2930, rule_2931, rule_2932, rule_2933, rule_2934, rule_2935, rule_2936, rule_2937, rule_2938, rule_2939, rule_2940, rule_2941, rule_2942, rule_2943, rule_2944, rule_2945, rule_2946, rule_2947, rule_2948, rule_2949, rule_2950, rule_2951, rule_2952, rule_2953, rule_2954, rule_2955, rule_2956, rule_2957, rule_2958, rule_2959, rule_2960, rule_2961, rule_2962, rule_2963, rule_2964, rule_2965, rule_2966, rule_2967, rule_2968, rule_2969, rule_2970, rule_2971, rule_2972, rule_2973, rule_2974, rule_2975, rule_2976, rule_2977, rule_2978, rule_2979, rule_2980, rule_2981, rule_2982, rule_2983, rule_2984, rule_2985, rule_2986, rule_2987, rule_2988, rule_2989, rule_2990, rule_2991, rule_2992, rule_2993, rule_2994, rule_2995, rule_2996, rule_2997, rule_2998, rule_2999, rule_3000, rule_3001, rule_3002, rule_3003, rule_3004, rule_3005, rule_3006, rule_3007, rule_3008, rule_3009, rule_3010, rule_3011, rule_3012, rule_3013, rule_3014, rule_3015, rule_3016, rule_3017, rule_3018, rule_3019, rule_3020, rule_3021, rule_3022, rule_3023, rule_3024, rule_3025, rule_3026, rule_3027, rule_3028, rule_3029, rule_3030, rule_3031, rule_3032, rule_3033, rule_3034, rule_3035, rule_3036, rule_3037, rule_3038, rule_3039, rule_3040, rule_3041, rule_3042, rule_3043, rule_3044, rule_3045, rule_3046, rule_3047, rule_3048, rule_3049, rule_3050, rule_3051, rule_3052, rule_3053, rule_3054, rule_3055, rule_3056, rule_3057, rule_3058, rule_3059, rule_3060, rule_3061, rule_3062, rule_3063, rule_3064, rule_3065, rule_3066, rule_3067, rule_3068, rule_3069, rule_3070, rule_3071, rule_3072, rule_3073, rule_3074, rule_3075, rule_3076, rule_3077, rule_3078, rule_3079, rule_3080, rule_3081, rule_3082, rule_3083, rule_3084, rule_3085, rule_3086, rule_3087, rule_3088, rule_3089, rule_3090, rule_3091, rule_3092, rule_3093, rule_3094, rule_3095, rule_3096, rule_3097, rule_3098, rule_3099, rule_3100, rule_3101, rule_3102, rule_3103, rule_3104, rule_3105, rule_3106, rule_3107, rule_3108, rule_3109, rule_3110, rule_3111, rule_3112, rule_3113, rule_3114, rule_3115, rule_3116, rule_3117, rule_3118, rule_3119, rule_3120, rule_3121, rule_3122, rule_3123, rule_3124, rule_3125, rule_3126, rule_3127, rule_3128, rule_3129, rule_3130, rule_3131, rule_3132, rule_3133, rule_3134, rule_3135, rule_3136, rule_3137, rule_3138, rule_3139, rule_3140, rule_3141, rule_3142, rule_3143, rule_3144, rule_3145, rule_3146, rule_3147, rule_3148, rule_3149, rule_3150, rule_3151, rule_3152, rule_3153, rule_3154, rule_3155, rule_3156, rule_3157, rule_3158, rule_3159, rule_3160, rule_3161, rule_3162, rule_3163, rule_3164, rule_3165, rule_3166, rule_3167, rule_3168, rule_3169, rule_3170, rule_3171, rule_3172, rule_3173, rule_3174, rule_3175, rule_3176, rule_3177, rule_3178, rule_3179, rule_3180, rule_3181, rule_3182, rule_3183, rule_3184, rule_3185, rule_3186, rule_3187, rule_3188, rule_3189, rule_3190, rule_3191, rule_3192, rule_3193, rule_3194, rule_3195, rule_3196, rule_3197, rule_3198, rule_3199, rule_3200, rule_3201, rule_3202, rule_3203, rule_3204, rule_3205, rule_3206, rule_3207, rule_3208, rule_3209, rule_3210, rule_3211, rule_3212, rule_3213, rule_3214, rule_3215, rule_3216, rule_3217, rule_3218, rule_3219, rule_3220, rule_3221, rule_3222, rule_3223, rule_3224, rule_3225, rule_3226, rule_3227, rule_3228, rule_3229, rule_3230, rule_3231, rule_3232, rule_3233, rule_3234, rule_3235, rule_3236, rule_3237, rule_3238, rule_3239, rule_3240, rule_3241, rule_3242, rule_3243, rule_3244, rule_3245, rule_3246, rule_3247, rule_3248, rule_3249, rule_3250, rule_3251, rule_3252, rule_3253, rule_3254, rule_3255, rule_3256, rule_3257, rule_3258, rule_3259, rule_3260, rule_3261, rule_3262, rule_3263, rule_3264, rule_3265, rule_3266, rule_3267, rule_3268, rule_3269, rule_3270, rule_3271, rule_3272, rule_3273, rule_3274, rule_3275, rule_3276, rule_3277, rule_3278, rule_3279, rule_3280, rule_3281, rule_3282, rule_3283, rule_3284, rule_3285, rule_3286, rule_3287, rule_3288, rule_3289, rule_3290, rule_3291, rule_3292, rule_3293, rule_3294, rule_3295, rule_3296, rule_3297, rule_3298, rule_3299, rule_3300, rule_3301, rule_3302, rule_3303, rule_3304, rule_3305, rule_3306, rule_3307, rule_3308, rule_3309, rule_3310, rule_3311, rule_3312, rule_3313, rule_3314, rule_3315, rule_3316, rule_3317, rule_3318, rule_3319, rule_3320, rule_3321, rule_3322, rule_3323, rule_3324, rule_3325, rule_3326, rule_3327, rule_3328, rule_3329, rule_3330, rule_3331, rule_3332, rule_3333, rule_3334, rule_3335, rule_3336, rule_3337, rule_3338, rule_3339, rule_3340, rule_3341, rule_3342, rule_3343, rule_3344, rule_3345, rule_3346, rule_3347, rule_3348, rule_3349, rule_3350, rule_3351, rule_3352, rule_3353, rule_3354, rule_3355, rule_3356, rule_3357, rule_3358, rule_3359, rule_3360, rule_3361, rule_3362, rule_3363, rule_3364, rule_3365, rule_3366, rule_3367, rule_3368, rule_3369, rule_3370, rule_3371, rule_3372, rule_3373, rule_3374, rule_3375, rule_3376, rule_3377, rule_3378, rule_3379, rule_3380, rule_3381, rule_3382, rule_3383, rule_3384, rule_3385, rule_3386, rule_3387, rule_3388, rule_3389, rule_3390, rule_3391, rule_3392, rule_3393, rule_3394, rule_3395, rule_3396, rule_3397, rule_3398, rule_3399, rule_3400, rule_3401, rule_3402, rule_3403, rule_3404, rule_3405, rule_3406, rule_3407, rule_3408, rule_3409, rule_3410, rule_3411, rule_3412, rule_3413, rule_3414, rule_3415, rule_3416, rule_3417, rule_3418, rule_3419, rule_3420, rule_3421, rule_3422, rule_3423, rule_3424, rule_3425, rule_3426, rule_3427, rule_3428, rule_3429, rule_3430, rule_3431, rule_3432, rule_3433, rule_3434, rule_3435, rule_3436, rule_3437, rule_3438, rule_3439, rule_3440, rule_3441, rule_3442, rule_3443, rule_3444, rule_3445, rule_3446, rule_3447, rule_3448, rule_3449, rule_3450, rule_3451, rule_3452, rule_3453, rule_3454, rule_3455, rule_3456, rule_3457, rule_3458, rule_3459, rule_3460, rule_3461, rule_3462, rule_3463, rule_3464, rule_3465, rule_3466, rule_3467, rule_3468, rule_3469, rule_3470, rule_3471, rule_3472, rule_3473, rule_3474, rule_3475, rule_3476, rule_3477, rule_3478, rule_3479, rule_3480, rule_3481, rule_3482, rule_3483, rule_3484, rule_3485, rule_3486, rule_3487, rule_3488, rule_3489, rule_3490, rule_3491, rule_3492, rule_3493, rule_3494, rule_3495, rule_3496, rule_3497, rule_3498, rule_3499, rule_3500, rule_3501, rule_3502, rule_3503, rule_3504, rule_3505, rule_3506, rule_3507, rule_3508, rule_3509, rule_3510, rule_3511, rule_3512, rule_3513, rule_3514, rule_3515, rule_3516, rule_3517, rule_3518, rule_3519, rule_3520, rule_3521, rule_3522, rule_3523, rule_3524, rule_3525, rule_3526, rule_3527, rule_3528, rule_3529, rule_3530, rule_3531, rule_3532, rule_3533, rule_3534, rule_3535, rule_3536, rule_3537, rule_3538, rule_3539, rule_3540, rule_3541, rule_3542, rule_3543, rule_3544, rule_3545, rule_3546, rule_3547, rule_3548, rule_3549, rule_3550, rule_3551, rule_3552, rule_3553, rule_3554, rule_3555, rule_3556, rule_3557, rule_3558, rule_3559, rule_3560, rule_3561, rule_3562, rule_3563, rule_3564, rule_3565, rule_3566, rule_3567, rule_3568, rule_3569, rule_3570, rule_3571, rule_3572, rule_3573, rule_3574, rule_3575, rule_3576, rule_3577, rule_3578, rule_3579, rule_3580, rule_3581, rule_3582, rule_3583, rule_3584, rule_3585, rule_3586, rule_3587, rule_3588, rule_3589, rule_3590, rule_3591, rule_3592, rule_3593, rule_3594, rule_3595, rule_3596, rule_3597, rule_3598, rule_3599, rule_3600, rule_3601, rule_3602, rule_3603, rule_3604, rule_3605, rule_3606, rule_3607, rule_3608, rule_3609, rule_3610, rule_3611, rule_3612, rule_3613, rule_3614, rule_3615, rule_3616, rule_3617, rule_3618, rule_3619, rule_3620, rule_3621, rule_3622, rule_3623, rule_3624, rule_3625, rule_3626, rule_3627, rule_3628, rule_3629, rule_3630, rule_3631, rule_3632, rule_3633, rule_3634, rule_3635, rule_3636, rule_3637, rule_3638, rule_3639, rule_3640, rule_3641, rule_3642, rule_3643, rule_3644, rule_3645, rule_3646, rule_3647, rule_3648, rule_3649, rule_3650, rule_3651, rule_3652, rule_3653, rule_3654, rule_3655, rule_3656, rule_3657, rule_3658, rule_3659, rule_3660, rule_3661, rule_3662, rule_3663, rule_3664, rule_3665, rule_3666, rule_3667, rule_3668, rule_3669, rule_3670, rule_3671, rule_3672, rule_3673, rule_3674, rule_3675, rule_3676, rule_3677, rule_3678, rule_3679, rule_3680, rule_3681, rule_3682, rule_3683, rule_3684, rule_3685, rule_3686, rule_3687, rule_3688, rule_3689, rule_3690, rule_3691, rule_3692, rule_3693, rule_3694, rule_3695, rule_3696, rule_3697, rule_3698, rule_3699, rule_3700, rule_3701, rule_3702, rule_3703, rule_3704, rule_3705, rule_3706, rule_3707, rule_3708, rule_3709, rule_3710, rule_3711, rule_3712, rule_3713, rule_3714, rule_3715, rule_3716, rule_3717, rule_3718, rule_3719, rule_3720, rule_3721, rule_3722, rule_3723, rule_3724, rule_3725, rule_3726, rule_3727, rule_3728, rule_3729, rule_3730, rule_3731, rule_3732, rule_3733, rule_3734, rule_3735, rule_3736, rule_3737, rule_3738, rule_3739, rule_3740, rule_3741, rule_3742, rule_3743, rule_3744, rule_3745, rule_3746, rule_3747, rule_3748, rule_3749, rule_3750, rule_3751, rule_3752, rule_3753, rule_3754, rule_3755, rule_3756, rule_3757, rule_3758, rule_3759, rule_3760, rule_3761, rule_3762, rule_3763, rule_3764, rule_3765, rule_3766, rule_3767, rule_3768, rule_3769, rule_3770, rule_3771, rule_3772, rule_3773, rule_3774, rule_3775, rule_3776, rule_3777, rule_3778, rule_3779, rule_3780, rule_3781, rule_3782, rule_3783, rule_3784, rule_3785, rule_3786, rule_3787, rule_3788, rule_3789, rule_3790, rule_3791, rule_3792, rule_3793, rule_3794, rule_3795, rule_3796, rule_3797, rule_3798, rule_3799, rule_3800, rule_3801, rule_3802, rule_3803, rule_3804, rule_3805, rule_3806, rule_3807, rule_3808, rule_3809, rule_3810, rule_3811, rule_3812, rule_3813, rule_3814, rule_3815, rule_3816, rule_3817, rule_3818, rule_3819, rule_3820, rule_3821, rule_3822, rule_3823, rule_3824, rule_3825, rule_3826, rule_3827, rule_3828, rule_3829, rule_3830, rule_3831, rule_3832, rule_3833, rule_3834, rule_3835, rule_3836, rule_3837, rule_3838, rule_3839, rule_3840, rule_3841, rule_3842, rule_3843, rule_3844, rule_3845, rule_3846, rule_3847, rule_3848, rule_3849, rule_3850, rule_3851, rule_3852, rule_3853, rule_3854, rule_3855, rule_3856, rule_3857, rule_3858, rule_3859, rule_3860, rule_3861, rule_3862, rule_3863, rule_3864, rule_3865, rule_3866, rule_3867, rule_3868, rule_3869, rule_3870, rule_3871, rule_3872, rule_3873, rule_3874, rule_3875, rule_3876, rule_3877, rule_3878, rule_3879, rule_3880, rule_3881, rule_3882, rule_3883, rule_3884, rule_3885, rule_3886, rule_3887, rule_3888, rule_3889, rule_3890, rule_3891, rule_3892, rule_3893, rule_3894, rule_3895, rule_3896, rule_3897, rule_3898, rule_3899, rule_3900, rule_3901, rule_3902, rule_3903, rule_3904, rule_3905, rule_3906, rule_3907, rule_3908, rule_3909, rule_3910, rule_3911, rule_3912, rule_3913, rule_3914, rule_3915, rule_3916, rule_3917, rule_3918, rule_3919, rule_3920, rule_3921, rule_3922, rule_3923, rule_3924, rule_3925, rule_3926, rule_3927, rule_3928, rule_3929, rule_3930, rule_3931, rule_3932, rule_3933, rule_3934, rule_3935, rule_3936, rule_3937, rule_3938, rule_3939, rule_3940, rule_3941, rule_3942, rule_3943, rule_3944, rule_3945, rule_3946, rule_3947, rule_3948, rule_3949, rule_3950, rule_3951, rule_3952, rule_3953, rule_3954, rule_3955, rule_3956, rule_3957, rule_3958, rule_3959, rule_3960, rule_3961, rule_3962, rule_3963, rule_3964, rule_3965, rule_3966, rule_3967, rule_3968, rule_3969, rule_3970, rule_3971, rule_3972, rule_3973, rule_3974, rule_3975, rule_3976, rule_3977, rule_3978, rule_3979, rule_3980, rule_3981, rule_3982, rule_3983, rule_3984, rule_3985, rule_3986, rule_3987, rule_3988, rule_3989, rule_3990, rule_3991, rule_3992, rule_3993, rule_3994, rule_3995, rule_3996, rule_3997, rule_3998, rule_3999, rule_4000, rule_4001, rule_4002, rule_4003, rule_4004, rule_4005, rule_4006, rule_4007, rule_4008, rule_4009, rule_4010, rule_4011, rule_4012, rule_4013, rule_4014, rule_4015, rule_4016, rule_4017, rule_4018, rule_4019, rule_4020, rule_4021, rule_4022, rule_4023, rule_4024, rule_4025, rule_4026, rule_4027, rule_4028, rule_4029, rule_4030, rule_4031, rule_4032, rule_4033, rule_4034, rule_4035, rule_4036, rule_4037, rule_4038, rule_4039, rule_4040, rule_4041, rule_4042, rule_4043, rule_4044, rule_4045, rule_4046, rule_4047, rule_4048, rule_4049, rule_4050, rule_4051, rule_4052, rule_4053, rule_4054, rule_4055, rule_4056, rule_4057, rule_4058, rule_4059, rule_4060, rule_4061, rule_4062, rule_4063, rule_4064, rule_4065, rule_4066, rule_4067, rule_4068, rule_4069, rule_4070, rule_4071, rule_4072, rule_4073, rule_4074, rule_4075, rule_4076, rule_4077, rule_4078, rule_4079, rule_4080, rule_4081, rule_4082, rule_4083, rule_4084, rule_4085, rule_4086, rule_4087, rule_4088, rule_4089, rule_4090, rule_4091, rule_4092, rule_4093, rule_4094, rule_4095, rule_4096, rule_4097, rule_4098, rule_4099, rule_4100, rule_4101, rule_4102, rule_4103, rule_4104, rule_4105, rule_4106, rule_4107, rule_4108, rule_4109, rule_4110, rule_4111, rule_4112, rule_4113, rule_4114, rule_4115, rule_4116, rule_4117, rule_4118, rule_4119, rule_4120, rule_4121, rule_4122, rule_4123, rule_4124, rule_4125, rule_4126, rule_4127, rule_4128, rule_4129, rule_4130, rule_4131, rule_4132, rule_4133, rule_4134, rule_4135, rule_4136, rule_4137, rule_4138, rule_4139, rule_4140, rule_4141, rule_4142, rule_4143, rule_4144, rule_4145, rule_4146, rule_4147, rule_4148, rule_4149, rule_4150, rule_4151, rule_4152, rule_4153, rule_4154, rule_4155, rule_4156, rule_4157, rule_4158, rule_4159, rule_4160, rule_4161, rule_4162, rule_4163, rule_4164, rule_4165, rule_4166, rule_4167, rule_4168, rule_4169, rule_4170, rule_4171, rule_4172, rule_4173, rule_4174, rule_4175, rule_4176, rule_4177, rule_4178, rule_4179, rule_4180, rule_4181, rule_4182, rule_4183, rule_4184, rule_4185, rule_4186, rule_4187, rule_4188, rule_4189, rule_4190, rule_4191, rule_4192, rule_4193, rule_4194, rule_4195, rule_4196, rule_4197, rule_4198, rule_4199, rule_4200, rule_4201, rule_4202, rule_4203, rule_4204, rule_4205, rule_4206, rule_4207, rule_4208, rule_4209, rule_4210, rule_4211, rule_4212, rule_4213, rule_4214, rule_4215, rule_4216, rule_4217, rule_4218, rule_4219, rule_4220, rule_4221, rule_4222, rule_4223, rule_4224, rule_4225, rule_4226, rule_4227, rule_4228, rule_4229, rule_4230, rule_4231, rule_4232, rule_4233, rule_4234, rule_4235, rule_4236, rule_4237, rule_4238, rule_4239, rule_4240, rule_4241, rule_4242, rule_4243, rule_4244, rule_4245, rule_4246, rule_4247, rule_4248, rule_4249, rule_4250, rule_4251, rule_4252, rule_4253, rule_4254, rule_4255, rule_4256, rule_4257, rule_4258, rule_4259, rule_4260, rule_4261, rule_4262, rule_4263, rule_4264, rule_4265, rule_4266, rule_4267, rule_4268, rule_4269, rule_4270, rule_4271, rule_4272, rule_4273, rule_4274, rule_4275, rule_4276, rule_4277, rule_4278, rule_4279, rule_4280, rule_4281, rule_4282, rule_4283, rule_4284, rule_4285, rule_4286, rule_4287, rule_4288, rule_4289, rule_4290, rule_4291, rule_4292, rule_4293, rule_4294, rule_4295, rule_4296, rule_4297, rule_4298, rule_4299, rule_4300, rule_4301, rule_4302, rule_4303, rule_4304, rule_4305, rule_4306, rule_4307, rule_4308, rule_4309, rule_4310, rule_4311, rule_4312, rule_4313, rule_4314, rule_4315, rule_4316, rule_4317, rule_4318, rule_4319, rule_4320, rule_4321, rule_4322, rule_4323, rule_4324, rule_4325, rule_4326, rule_4327, rule_4328, rule_4329, rule_4330, rule_4331, rule_4332, rule_4333, rule_4334, rule_4335, rule_4336, rule_4337, rule_4338, rule_4339, rule_4340, rule_4341, rule_4342, rule_4343, rule_4344, rule_4345, rule_4346, rule_4347, rule_4348, rule_4349, rule_4350, rule_4351, rule_4352, rule_4353, rule_4354, rule_4355, rule_4356, rule_4357, rule_4358, rule_4359, rule_4360, rule_4361, rule_4362, rule_4363, rule_4364, rule_4365, rule_4366, rule_4367, rule_4368, rule_4369, rule_4370, rule_4371, rule_4372, rule_4373, rule_4374, rule_4375, rule_4376, rule_4377, rule_4378, rule_4379, rule_4380, rule_4381, rule_4382, rule_4383, rule_4384, rule_4385, rule_4386, rule_4387, rule_4388, rule_4389, rule_4390, rule_4391, rule_4392, rule_4393, rule_4394, rule_4395, rule_4396, rule_4397, rule_4398, rule_4399, rule_4400, rule_4401, rule_4402, rule_4403, rule_4404, rule_4405, rule_4406, rule_4407, rule_4408, rule_4409, rule_4410, rule_4411, rule_4412, rule_4413, rule_4414, rule_4415, rule_4416, rule_4417, rule_4418, rule_4419, rule_4420, rule_4421, rule_4422, rule_4423, rule_4424, rule_4425, rule_4426, rule_4427, rule_4428, rule_4429, rule_4430, rule_4431, rule_4432, rule_4433, rule_4434, rule_4435, rule_4436, rule_4437, rule_4438, rule_4439, rule_4440, rule_4441, rule_4442, rule_4443, rule_4444, rule_4445, rule_4446, rule_4447, rule_4448, rule_4449, rule_4450, rule_4451, rule_4452, rule_4453, rule_4454, rule_4455, rule_4456, rule_4457, rule_4458, rule_4459, rule_4460, rule_4461, rule_4462, rule_4463, rule_4464, rule_4465, rule_4466, rule_4467, rule_4468, rule_4469, rule_4470, rule_4471, rule_4472, rule_4473, rule_4474, rule_4475, rule_4476, rule_4477, rule_4478, rule_4479, rule_4480, rule_4481, rule_4482, rule_4483, rule_4484, rule_4485, rule_4486, rule_4487, rule_4488, rule_4489, rule_4490, rule_4491, rule_4492, rule_4493, rule_4494, rule_4495, rule_4496, rule_4497, rule_4498, rule_4499, rule_4500, rule_4501, rule_4502, rule_4503, rule_4504, rule_4505, rule_4506, rule_4507, rule_4508, rule_4509, rule_4510, rule_4511, rule_4512, rule_4513, rule_4514, rule_4515, rule_4516, rule_4517, rule_4518, rule_4519, rule_4520, rule_4521, rule_4522, rule_4523, rule_4524, rule_4525, rule_4526, rule_4527, rule_4528, rule_4529, rule_4530, rule_4531, rule_4532, rule_4533, rule_4534, rule_4535, rule_4536, rule_4537, rule_4538, rule_4539, rule_4540, rule_4541, rule_4542, rule_4543, rule_4544, rule_4545, rule_4546, rule_4547, rule_4548, rule_4549, rule_4550, rule_4551, rule_4552, rule_4553, rule_4554, rule_4555, rule_4556, rule_4557, rule_4558, rule_4559, rule_4560, rule_4561, rule_4562, rule_4563, rule_4564, rule_4565, rule_4566, rule_4567, rule_4568, rule_4569, rule_4570, rule_4571, rule_4572, rule_4573, rule_4574, rule_4575, rule_4576, rule_4577, rule_4578, rule_4579, rule_4580, rule_4581, rule_4582, rule_4583, rule_4584, rule_4585, rule_4586, rule_4587, rule_4588, rule_4589, rule_4590, rule_4591, rule_4592, rule_4593, rule_4594, rule_4595, rule_4596, rule_4597, rule_4598, rule_4599, rule_4600, rule_4601, rule_4602, rule_4603, rule_4604, rule_4605, rule_4606, rule_4607, rule_4608, rule_4609, rule_4610, rule_4611, rule_4612, rule_4613, rule_4614, rule_4615, rule_4616, rule_4617, rule_4618, rule_4619, rule_4620, rule_4621, rule_4622, rule_4623, rule_4624, rule_4625, rule_4626, rule_4627, rule_4628, rule_4629, rule_4630, rule_4631, rule_4632, rule_4633, rule_4634, rule_4635, rule_4636, rule_4637, rule_4638, rule_4639, rule_4640, rule_4641, rule_4642, rule_4643, rule_4644, rule_4645, rule_4646, rule_4647, rule_4648, rule_4649, rule_4650, rule_4651, rule_4652, rule_4653, rule_4654, rule_4655, rule_4656, rule_4657, rule_4658, rule_4659, rule_4660, rule_4661, rule_4662, rule_4663, rule_4664, rule_4665, rule_4666, rule_4667, rule_4668, rule_4669, rule_4670, rule_4671, rule_4672, rule_4673, rule_4674, rule_4675, rule_4676, rule_4677, rule_4678, rule_4679, rule_4680, rule_4681, rule_4682, rule_4683, rule_4684, rule_4685, rule_4686, rule_4687, rule_4688, rule_4689, rule_4690, rule_4691, rule_4692, rule_4693, rule_4694, rule_4695, rule_4696, rule_4697, rule_4698, rule_4699, rule_4700, rule_4701, rule_4702, rule_4703, rule_4704, rule_4705, rule_4706, rule_4707, rule_4708, rule_4709, rule_4710, rule_4711, rule_4712, rule_4713, rule_4714, rule_4715, rule_4716, rule_4717, rule_4718, rule_4719, rule_4720, rule_4721, rule_4722, rule_4723, rule_4724, rule_4725, rule_4726, rule_4727, rule_4728, rule_4729, rule_4730, rule_4731, rule_4732, rule_4733, rule_4734, rule_4735, rule_4736, rule_4737, rule_4738, rule_4739, rule_4740, rule_4741, rule_4742, rule_4743, rule_4744, rule_4745, rule_4746, rule_4747, rule_4748, rule_4749, rule_4750, rule_4751, rule_4752, rule_4753, rule_4754, rule_4755, rule_4756, rule_4757, rule_4758, rule_4759, rule_4760, rule_4761, rule_4762, rule_4763, rule_4764, rule_4765, rule_4766, rule_4767, rule_4768, rule_4769, rule_4770, rule_4771, rule_4772, rule_4773, rule_4774, rule_4775, rule_4776, rule_4777, rule_4778, rule_4779, rule_4780, rule_4781, rule_4782, rule_4783, rule_4784, rule_4785, rule_4786, rule_4787, rule_4788, rule_4789, rule_4790, rule_4791, rule_4792, rule_4793, rule_4794, rule_4795, rule_4796, rule_4797, rule_4798, rule_4799, rule_4800, rule_4801, rule_4802, rule_4803, rule_4804, rule_4805, rule_4806, rule_4807, rule_4808, rule_4809, rule_4810, rule_4811, rule_4812, rule_4813, rule_4814, rule_4815, rule_4816, rule_4817, rule_4818, rule_4819, rule_4820, rule_4821, rule_4822, rule_4823, rule_4824, rule_4825, rule_4826, rule_4827, rule_4828, rule_4829, rule_4830, rule_4831, rule_4832, rule_4833, rule_4834, rule_4835, rule_4836, rule_4837, rule_4838, rule_4839, rule_4840, rule_4841, rule_4842, rule_4843, rule_4844, rule_4845, rule_4846, rule_4847, rule_4848, rule_4849, rule_4850, rule_4851, rule_4852, rule_4853, rule_4854, rule_4855, rule_4856, rule_4857, rule_4858, rule_4859, rule_4860, rule_4861, rule_4862, rule_4863, rule_4864, rule_4865, rule_4866, rule_4867, rule_4868, rule_4869, rule_4870, rule_4871, rule_4872, rule_4873, rule_4874, rule_4875, rule_4876, rule_4877, rule_4878, rule_4879, rule_4880, rule_4881, rule_4882, rule_4883, rule_4884, rule_4885, rule_4886, rule_4887, rule_4888, rule_4889, rule_4890, rule_4891, rule_4892, rule_4893, rule_4894, rule_4895, rule_4896, rule_4897, rule_4898, rule_4899, rule_4900, rule_4901, rule_4902, rule_4903, rule_4904, rule_4905, rule_4906, rule_4907, rule_4908, rule_4909, rule_4910, rule_4911, rule_4912, rule_4913, rule_4914, rule_4915, rule_4916, rule_4917, rule_4918, rule_4919, rule_4920, rule_4921, rule_4922, rule_4923, rule_4924, rule_4925, rule_4926, rule_4927, rule_4928, rule_4929, rule_4930, rule_4931, rule_4932, rule_4933, rule_4934, rule_4935, rule_4936, rule_4937, rule_4938, rule_4939, rule_4940, rule_4941, rule_4942, rule_4943, rule_4944, rule_4945, rule_4946, rule_4947, rule_4948, rule_4949, rule_4950, rule_4951, rule_4952, rule_4953, rule_4954, rule_4955, rule_4956, rule_4957, rule_4958, rule_4959, rule_4960, rule_4961, rule_4962, rule_4963, rule_4964, rule_4965, rule_4966, rule_4967, rule_4968, rule_4969, rule_4970, rule_4971, rule_4972, rule_4973, rule_4974, rule_4975, rule_4976, rule_4977, rule_4978, rule_4979, rule_4980, rule_4981, rule_4982, rule_4983, rule_4984, rule_4985, rule_4986, rule_4987, rule_4988, rule_4989, rule_4990, rule_4991, rule_4992, rule_4993, rule_4994, rule_4995, rule_4996, rule_4997, rule_4998, rule_4999, rule_5000, rule_5001, rule_5002, rule_5003, rule_5004, rule_5005, rule_5006, rule_5007, rule_5008, rule_5009, rule_5010, rule_5011, rule_5012, rule_5013, rule_5014, rule_5015, rule_5016, rule_5017, rule_5018, rule_5019, rule_5020, rule_5021, rule_5022, rule_5023, rule_5024, rule_5025, rule_5026, rule_5027, rule_5028, rule_5029, rule_5030, rule_5031, rule_5032, rule_5033, rule_5034, rule_5035, rule_5036, rule_5037, rule_5038, rule_5039, rule_5040, rule_5041, rule_5042, rule_5043, rule_5044, rule_5045, rule_5046, rule_5047, rule_5048, rule_5049, rule_5050, rule_5051, rule_5052, rule_5053, rule_5054, rule_5055, rule_5056, rule_5057, rule_5058, rule_5059, rule_5060, rule_5061, rule_5062, rule_5063, rule_5064, rule_5065, rule_5066, rule_5067, rule_5068, rule_5069, rule_5070, rule_5071, rule_5072, rule_5073, rule_5074, rule_5075, rule_5076, rule_5077, rule_5078, rule_5079, rule_5080, rule_5081, rule_5082, rule_5083, rule_5084, rule_5085, rule_5086, rule_5087, rule_5088, rule_5089, rule_5090, rule_5091, rule_5092, rule_5093, rule_5094, rule_5095, rule_5096, rule_5097, rule_5098, rule_5099, rule_5100, rule_5101, rule_5102, rule_5103, rule_5104, rule_5105, rule_5106, rule_5107, rule_5108, rule_5109, rule_5110, rule_5111, rule_5112, rule_5113, rule_5114, rule_5115, rule_5116, rule_5117, rule_5118, rule_5119, rule_5120, rule_5121, rule_5122, rule_5123, rule_5124, rule_5125, rule_5126, rule_5127, rule_5128, rule_5129, rule_5130, rule_5131, rule_5132, rule_5133, rule_5134, rule_5135, rule_5136, rule_5137, rule_5138, rule_5139, rule_5140, rule_5141, rule_5142, rule_5143, rule_5144, rule_5145, rule_5146, rule_5147, rule_5148, rule_5149, rule_5150, rule_5151, rule_5152, rule_5153, rule_5154, rule_5155, rule_5156, rule_5157, rule_5158, rule_5159, rule_5160, rule_5161, rule_5162, rule_5163, rule_5164, rule_5165, rule_5166, rule_5167, rule_5168, rule_5169, rule_5170, rule_5171, rule_5172, rule_5173, rule_5174, rule_5175, rule_5176, rule_5177, rule_5178, rule_5179, rule_5180, rule_5181, rule_5182, rule_5183, rule_5184, rule_5185, rule_5186, rule_5187, rule_5188, rule_5189, rule_5190, rule_5191, rule_5192, rule_5193, rule_5194, rule_5195, rule_5196, rule_5197, rule_5198, rule_5199, rule_5200, rule_5201, rule_5202, rule_5203, rule_5204, rule_5205, rule_5206, rule_5207, rule_5208, rule_5209, rule_5210, rule_5211, rule_5212, rule_5213, rule_5214, rule_5215, rule_5216, rule_5217, rule_5218, rule_5219, rule_5220, rule_5221, rule_5222, rule_5223, rule_5224, rule_5225, rule_5226, rule_5227, rule_5228, rule_5229, rule_5230, rule_5231, rule_5232, rule_5233, rule_5234, rule_5235, rule_5236, rule_5237, rule_5238, rule_5239, rule_5240, rule_5241, rule_5242, rule_5243, rule_5244, rule_5245, rule_5246, rule_5247, rule_5248, rule_5249, rule_5250, rule_5251, rule_5252, rule_5253, rule_5254, rule_5255, rule_5256, rule_5257, rule_5258, rule_5259, rule_5260, rule_5261, rule_5262, rule_5263, rule_5264, rule_5265, rule_5266, rule_5267, rule_5268, rule_5269, rule_5270, rule_5271, rule_5272, rule_5273, rule_5274, rule_5275, rule_5276, rule_5277, rule_5278, rule_5279, rule_5280, rule_5281, rule_5282, rule_5283, rule_5284, rule_5285, rule_5286, rule_5287, rule_5288, rule_5289, rule_5290, rule_5291, rule_5292, rule_5293, rule_5294, rule_5295, rule_5296, rule_5297, rule_5298, rule_5299, rule_5300, rule_5301, rule_5302, rule_5303, rule_5304, rule_5305, rule_5306, rule_5307, rule_5308, rule_5309, rule_5310, rule_5311, rule_5312, rule_5313, rule_5314, rule_5315, rule_5316, rule_5317, rule_5318, rule_5319, rule_5320, rule_5321, rule_5322, rule_5323, rule_5324, rule_5325, rule_5326, rule_5327, rule_5328, rule_5329, rule_5330, rule_5331, rule_5332, rule_5333, rule_5334, rule_5335, rule_5336, rule_5337, rule_5338, rule_5339, rule_5340, rule_5341, rule_5342, rule_5343, rule_5344, rule_5345, rule_5346, rule_5347, rule_5348, rule_5349, rule_5350, rule_5351, rule_5352, rule_5353, rule_5354, rule_5355, rule_5356, rule_5357, rule_5358, rule_5359, rule_5360, rule_5361, rule_5362, rule_5363, rule_5364, rule_5365, rule_5366, rule_5367, rule_5368, rule_5369, rule_5370, rule_5371, rule_5372, rule_5373, rule_5374, rule_5375, rule_5376, rule_5377, rule_5378, rule_5379, rule_5380, rule_5381, rule_5382, rule_5383, rule_5384, rule_5385, rule_5386, rule_5387, rule_5388, rule_5389, rule_5390, rule_5391, rule_5392, rule_5393, rule_5394, rule_5395, rule_5396, rule_5397, rule_5398, rule_5399, rule_5400, rule_5401, rule_5402, rule_5403, rule_5404, rule_5405, rule_5406, rule_5407, rule_5408, rule_5409, rule_5410, rule_5411, rule_5412, rule_5413, rule_5414, rule_5415, rule_5416, rule_5417, rule_5418, rule_5419, rule_5420, rule_5421, rule_5422, rule_5423, rule_5424, rule_5425, rule_5426, rule_5427, rule_5428, rule_5429, rule_5430, rule_5431, rule_5432, rule_5433, rule_5434, rule_5435, rule_5436, rule_5437, rule_5438, rule_5439, rule_5440, rule_5441, rule_5442, rule_5443, rule_5444, rule_5445, rule_5446, rule_5447, rule_5448, rule_5449, rule_5450, rule_5451, rule_5452, rule_5453, rule_5454, rule_5455, rule_5456, rule_5457, rule_5458, rule_5459, rule_5460, rule_5461, rule_5462, rule_5463, rule_5464, rule_5465, rule_5466, rule_5467, rule_5468, rule_5469, rule_5470, rule_5471, rule_5472, rule_5473, rule_5474, rule_5475, rule_5476, rule_5477, rule_5478, rule_5479, rule_5480, rule_5481, rule_5482, rule_5483, rule_5484, rule_5485, rule_5486, rule_5487, rule_5488, rule_5489, rule_5490, rule_5491, rule_5492, rule_5493, rule_5494, rule_5495, rule_5496, rule_5497, rule_5498, rule_5499, rule_5500, rule_5501, rule_5502, rule_5503, rule_5504, rule_5505, rule_5506, rule_5507, rule_5508, rule_5509, rule_5510, rule_5511, rule_5512, rule_5513, rule_5514, rule_5515, rule_5516, rule_5517, rule_5518, rule_5519, rule_5520, rule_5521, rule_5522, rule_5523, rule_5524, rule_5525, rule_5526, rule_5527, rule_5528, rule_5529, rule_5530, rule_5531, rule_5532, rule_5533, rule_5534, rule_5535, rule_5536, rule_5537, rule_5538, rule_5539, rule_5540, rule_5541, rule_5542, rule_5543, rule_5544, rule_5545, rule_5546, rule_5547, rule_5548, rule_5549, rule_5550, rule_5551, rule_5552, rule_5553, rule_5554, rule_5555, rule_5556, rule_5557, rule_5558, rule_5559, rule_5560, rule_5561, rule_5562, rule_5563, rule_5564, rule_5565, rule_5566, rule_5567, rule_5568, rule_5569, rule_5570, rule_5571, rule_5572, rule_5573, rule_5574, rule_5575, rule_5576, rule_5577, rule_5578, rule_5579, rule_5580, rule_5581, rule_5582, rule_5583, rule_5584, rule_5585, rule_5586, rule_5587, rule_5588, rule_5589, rule_5590, rule_5591, rule_5592, rule_5593, rule_5594, rule_5595, rule_5596, rule_5597, rule_5598, rule_5599, rule_5600, rule_5601, rule_5602, rule_5603, rule_5604, rule_5605, rule_5606, rule_5607, rule_5608, rule_5609, rule_5610, rule_5611, rule_5612, rule_5613, rule_5614, rule_5615, rule_5616, rule_5617, rule_5618, rule_5619, rule_5620, rule_5621, rule_5622, rule_5623, rule_5624, rule_5625, rule_5626, rule_5627, rule_5628, rule_5629, rule_5630, rule_5631, rule_5632, rule_5633, rule_5634, rule_5635, rule_5636, rule_5637, rule_5638, rule_5639, rule_5640, rule_5641, rule_5642, rule_5643, rule_5644, rule_5645, rule_5646, rule_5647, rule_5648, rule_5649, rule_5650, rule_5651, rule_5652, rule_5653, rule_5654, rule_5655, rule_5656, rule_5657, rule_5658, rule_5659, rule_5660, rule_5661, rule_5662, rule_5663, rule_5664, rule_5665, rule_5666, rule_5667, rule_5668, rule_5669, rule_5670, rule_5671, rule_5672, rule_5673, rule_5674, rule_5675, rule_5676, rule_5677, rule_5678, rule_5679, rule_5680, rule_5681, rule_5682, rule_5683, rule_5684, rule_5685, rule_5686, rule_5687, rule_5688, rule_5689, rule_5690, rule_5691, rule_5692, rule_5693, rule_5694, rule_5695, rule_5696, rule_5697, rule_5698, rule_5699, rule_5700, rule_5701, rule_5702, rule_5703, rule_5704, rule_5705, rule_5706, rule_5707, rule_5708, rule_5709, rule_5710, rule_5711, rule_5712, rule_5713, rule_5714, rule_5715, rule_5716, rule_5717, rule_5718, rule_5719, rule_5720, rule_5721, rule_5722, rule_5723, rule_5724, rule_5725, rule_5726, rule_5727, rule_5728, rule_5729, rule_5730, rule_5731, rule_5732, rule_5733, rule_5734, rule_5735, rule_5736, rule_5737, rule_5738, rule_5739, rule_5740, rule_5741, rule_5742, rule_5743, rule_5744, rule_5745, rule_5746, rule_5747, rule_5748, rule_5749, rule_5750, rule_5751, rule_5752, rule_5753, rule_5754, rule_5755, rule_5756, rule_5757, rule_5758, rule_5759, rule_5760, rule_5761, rule_5762, rule_5763, rule_5764, rule_5765, rule_5766, rule_5767, rule_5768, rule_5769, rule_5770, rule_5771, rule_5772, rule_5773, rule_5774, rule_5775, rule_5776, rule_5777, rule_5778, rule_5779, rule_5780, rule_5781, rule_5782, rule_5783, rule_5784, rule_5785, rule_5786, rule_5787, rule_5788, rule_5789, rule_5790, rule_5791, rule_5792, rule_5793, rule_5794, rule_5795, rule_5796, rule_5797, rule_5798, rule_5799, rule_5800, rule_5801, rule_5802, rule_5803, rule_5804, rule_5805, rule_5806, rule_5807, rule_5808, rule_5809, rule_5810, rule_5811, rule_5812, rule_5813, rule_5814, rule_5815, rule_5816, rule_5817, rule_5818, rule_5819, rule_5820, rule_5821, rule_5822, rule_5823, rule_5824, rule_5825, rule_5826, rule_5827, rule_5828, rule_5829, rule_5830, rule_5831, rule_5832, rule_5833, rule_5834, rule_5835, rule_5836, rule_5837, rule_5838, rule_5839, rule_5840, rule_5841, rule_5842, rule_5843, rule_5844, rule_5845, rule_5846, rule_5847, rule_5848, rule_5849, rule_5850, rule_5851, rule_5852, rule_5853, rule_5854, rule_5855, rule_5856, rule_5857, rule_5858, rule_5859, rule_5860, rule_5861, rule_5862, rule_5863, rule_5864, rule_5865, rule_5866, rule_5867, rule_5868, rule_5869, rule_5870, rule_5871, rule_5872, rule_5873, rule_5874, rule_5875, rule_5876, rule_5877, rule_5878, rule_5879, rule_5880, rule_5881, rule_5882, rule_5883, rule_5884, rule_5885, rule_5886, rule_5887, rule_5888, rule_5889, rule_5890, rule_5891, rule_5892, rule_5893, rule_5894, rule_5895, rule_5896, rule_5897, rule_5898, rule_5899, rule_5900, rule_5901, rule_5902, rule_5903, rule_5904, rule_5905, rule_5906, rule_5907, rule_5908, rule_5909, rule_5910, rule_5911, rule_5912, rule_5913, rule_5914, rule_5915, rule_5916, rule_5917, rule_5918, rule_5919, rule_5920, rule_5921, rule_5922, rule_5923, rule_5924, rule_5925, rule_5926, rule_5927, rule_5928, rule_5929, rule_5930, rule_5931, rule_5932, rule_5933, rule_5934, rule_5935, rule_5936, rule_5937, rule_5938, rule_5939, rule_5940, rule_5941, rule_5942, rule_5943, rule_5944, rule_5945, rule_5946, rule_5947, rule_5948, rule_5949, rule_5950, rule_5951, rule_5952, rule_5953, rule_5954, rule_5955, rule_5956, rule_5957, rule_5958, rule_5959, rule_5960, rule_5961, rule_5962, rule_5963, rule_5964, rule_5965, rule_5966, rule_5967, rule_5968, rule_5969, rule_5970, rule_5971, rule_5972, rule_5973, rule_5974, rule_5975, rule_5976, rule_5977, rule_5978, rule_5979, rule_5980, rule_5981, rule_5982, rule_5983, rule_5984, rule_5985, rule_5986, rule_5987, rule_5988, rule_5989, rule_5990, rule_5991, rule_5992, rule_5993, rule_5994, rule_5995, rule_5996, rule_5997, rule_5998, rule_5999, rule_6000, rule_6001, rule_6002, rule_6003, rule_6004, rule_6005, rule_6006, rule_6007, rule_6008, rule_6009, rule_6010, rule_6011, rule_6012, rule_6013, rule_6014, rule_6015, rule_6016, rule_6017, rule_6018, rule_6019, rule_6020, rule_6021, rule_6022, rule_6023, rule_6024, rule_6025, rule_6026, rule_6027, rule_6028, rule_6029, rule_6030, rule_6031, rule_6032, rule_6033, rule_6034, rule_6035, rule_6036, rule_6037, rule_6038, rule_6039, rule_6040, rule_6041, rule_6042, rule_6043, rule_6044, rule_6045, rule_6046, rule_6047, rule_6048, rule_6049, rule_6050, rule_6051, rule_6052, rule_6053, rule_6054, rule_6055, rule_6056, rule_6057, rule_6058, rule_6059, rule_6060, rule_6061, rule_6062, rule_6063, rule_6064, rule_6065, rule_6066, rule_6067, rule_6068, rule_6069, rule_6070, rule_6071, rule_6072, rule_6073, rule_6074, rule_6075, rule_6076, rule_6077, rule_6078, rule_6079, rule_6080, rule_6081, rule_6082, rule_6083, rule_6084, rule_6085, rule_6086, rule_6087, rule_6088, rule_6089, rule_6090, rule_6091, rule_6092, rule_6093, rule_6094, rule_6095, rule_6096, rule_6097, rule_6098, rule_6099, rule_6100, rule_6101, rule_6102, rule_6103, rule_6104, rule_6105, rule_6106, rule_6107, rule_6108, rule_6109, rule_6110, rule_6111, rule_6112, rule_6113, rule_6114, rule_6115, rule_6116, rule_6117, rule_6118, rule_6119, rule_6120, rule_6121, rule_6122, rule_6123, rule_6124, rule_6125, rule_6126, rule_6127, rule_6128, rule_6129, rule_6130, rule_6131, rule_6132, rule_6133, rule_6134, rule_6135, rule_6136, rule_6137, rule_6138, rule_6139, rule_6140, rule_6141, rule_6142, rule_6143, rule_6144, rule_6145, rule_6146, rule_6147, rule_6148, rule_6149, rule_6150, rule_6151, rule_6152, rule_6153, rule_6154, rule_6155, rule_6156, rule_6157, rule_6158, rule_6159, rule_6160, rule_6161, rule_6162, rule_6163, rule_6164, rule_6165, rule_6166, rule_6167, rule_6168, rule_6169, rule_6170, rule_6171, rule_6172, rule_6173, rule_6174, rule_6175, rule_6176, rule_6177, rule_6178, rule_6179, rule_6180, rule_6181, rule_6182, rule_6183, rule_6184, rule_6185, rule_6186, rule_6187, rule_6188, rule_6189, rule_6190, rule_6191, rule_6192, rule_6193, rule_6194, rule_6195, rule_6196, rule_6197, rule_6198, rule_6199, rule_6200, rule_6201, rule_6202, rule_6203, rule_6204, rule_6205, rule_6206, rule_6207, rule_6208, rule_6209, rule_6210, rule_6211, rule_6212, rule_6213, rule_6214, rule_6215, rule_6216, rule_6217, rule_6218, rule_6219, rule_6220, rule_6221, rule_6222, rule_6223, rule_6224, rule_6225, rule_6226, rule_6227, rule_6228, rule_6229, rule_6230, rule_6231, rule_6232, rule_6233, rule_6234, rule_6235, rule_6236, rule_6237, rule_6238, rule_6239, rule_6240, rule_6241, rule_6242, rule_6243, rule_6244, rule_6245, rule_6246, rule_6247, rule_6248, rule_6249, rule_6250, rule_6251, rule_6252, rule_6253, rule_6254, rule_6255, rule_6256, rule_6257, rule_6258, rule_6259, rule_6260, rule_6261, rule_6262, rule_6263, rule_6264, rule_6265, rule_6266, rule_6267, rule_6268, rule_6269, rule_6270, rule_6271, rule_6272, rule_6273, rule_6274, rule_6275, rule_6276, rule_6277, rule_6278, rule_6279, rule_6280, rule_6281, rule_6282, rule_6283, rule_6284, rule_6285, rule_6286, rule_6287, rule_6288, rule_6289, rule_6290, rule_6291, rule_6292, rule_6293, rule_6294, rule_6295, rule_6296, rule_6297, rule_6298, rule_6299, rule_6300, rule_6301, rule_6302, rule_6303, rule_6304, rule_6305, rule_6306, rule_6307, rule_6308, rule_6309, rule_6310, rule_6311, rule_6312, rule_6313, rule_6314, rule_6315, rule_6316, rule_6317, rule_6318, rule_6319, rule_6320, rule_6321, rule_6322, rule_6323, rule_6324, rule_6325, rule_6326, rule_6327, rule_6328, rule_6329, rule_6330, rule_6331, rule_6332, rule_6333, rule_6334, rule_6335, rule_6336, rule_6337, rule_6338, rule_6339, rule_6340, rule_6341, rule_6342, rule_6343, rule_6344, rule_6345, rule_6346, rule_6347, rule_6348, rule_6349, rule_6350, rule_6351, rule_6352, rule_6353, rule_6354, rule_6355, rule_6356, rule_6357, rule_6358, rule_6359, rule_6360, rule_6361, rule_6362, rule_6363, rule_6364, rule_6365, rule_6366, rule_6367, rule_6368, rule_6369, rule_6370, rule_6371, rule_6372, rule_6373, rule_6374, rule_6375, rule_6376, rule_6377, rule_6378, rule_6379, rule_6380, rule_6381, rule_6382, rule_6383, rule_6384, rule_6385, rule_6386, rule_6387, rule_6388, rule_6389, rule_6390, rule_6391, rule_6392, rule_6393, rule_6394, rule_6395, rule_6396, rule_6397, rule_6398, rule_6399, rule_6400, rule_6401, rule_6402, rule_6403, rule_6404, rule_6405, rule_6406, rule_6407, rule_6408, rule_6409, rule_6410, rule_6411, rule_6412, rule_6413, rule_6414, rule_6415, rule_6416, rule_6417, rule_6418, rule_6419, rule_6420, rule_6421, rule_6422, rule_6423, rule_6424, rule_6425, rule_6426, rule_6427, rule_6428, rule_6429, rule_6430, rule_6431, rule_6432, rule_6433, rule_6434, rule_6435, rule_6436, rule_6437, rule_6438, rule_6439, rule_6440, rule_6441, rule_6442, rule_6443, rule_6444, rule_6445, rule_6446, rule_6447, rule_6448, rule_6449, rule_6450, rule_6451, rule_6452, rule_6453, rule_6454, rule_6455, rule_6456, rule_6457, rule_6458, rule_6459, rule_6460, rule_6461, rule_6462, rule_6463, rule_6464, rule_6465, rule_6466, rule_6467, rule_6468, rule_6469, rule_6470, rule_6471, rule_6472, rule_6473, rule_6474, rule_6475, rule_6476, rule_6477, rule_6478, rule_6479, rule_6480, rule_6481, rule_6482, rule_6483, rule_6484, rule_6485, rule_6486, rule_6487, rule_6488, rule_6489, rule_6490, rule_6491, rule_6492, rule_6493, rule_6494, rule_6495, rule_6496, rule_6497, rule_6498, rule_6499, rule_6500, rule_6501, rule_6502, rule_6503, rule_6504, rule_6505, rule_6506, rule_6507, rule_6508, rule_6509, rule_6510, rule_6511, rule_6512, rule_6513, rule_6514, rule_6515, rule_6516, rule_6517, rule_6518, rule_6519, rule_6520, rule_6521, rule_6522, rule_6523, rule_6524, rule_6525, rule_6526, rule_6527, rule_6528, rule_6529, rule_6530, rule_6531, rule_6532, rule_6533, rule_6534, rule_6535, rule_6536, rule_6537, rule_6538, rule_6539, rule_6540, rule_6541, rule_6542, rule_6543, rule_6544, rule_6545, rule_6546, rule_6547, rule_6548, rule_6549, rule_6550, rule_6551, rule_6552, rule_6553, rule_6554, rule_6555, rule_6556, rule_6557, rule_6558, rule_6559, rule_6560, rule_6561, rule_6562, rule_6563, rule_6564, rule_6565, rule_6566, rule_6567, rule_6568, rule_6569, rule_6570, rule_6571, rule_6572, rule_6573, rule_6574, rule_6575, rule_6576, rule_6577, rule_6578, rule_6579, rule_6580, rule_6581, rule_6582, rule_6583, rule_6584, rule_6585, rule_6586, rule_6587, rule_6588, rule_6589, rule_6590, rule_6591, rule_6592, rule_6593, rule_6594, rule_6595, rule_6596, rule_6597, rule_6598, rule_6599, rule_6600, rule_6601, rule_6602, rule_6603, rule_6604, rule_6605, rule_6606, rule_6607, rule_6608, rule_6609, rule_6610, rule_6611, rule_6612, rule_6613, rule_6614, rule_6615, rule_6616, rule_6617, rule_6618, rule_6619, rule_6620, rule_6621, rule_6622, rule_6623, rule_6624, rule_6625, rule_6626, rule_6627, rule_6628, rule_6629, rule_6630, rule_6631, rule_6632, rule_6633, rule_6634, rule_6635, rule_6636, rule_6637, rule_6638, rule_6639, rule_6640, rule_6641, rule_6642, rule_6643, rule_6644, rule_6645, rule_6646, rule_6647, rule_6648, rule_6649, rule_6650, rule_6651, rule_6652, rule_6653, rule_6654, rule_6655, rule_6656, rule_6657, rule_6658, rule_6659, rule_6660, rule_6661, rule_6662, rule_6663, rule_6664, rule_6665, rule_6666, rule_6667, rule_6668, rule_6669, rule_6670, rule_6671, rule_6672, rule_6673, rule_6674, rule_6675, rule_6676, rule_6677, rule_6678, rule_6679, rule_6680, rule_6681, rule_6682, rule_6683, rule_6684, rule_6685, rule_6686, rule_6687, rule_6688, rule_6689, rule_6690, rule_6691, rule_6692, rule_6693, rule_6694, rule_6695, rule_6696, rule_6697, rule_6698, rule_6699, rule_6700, rule_6701, rule_6702, rule_6703, rule_6704, rule_6705, rule_6706, rule_6707, rule_6708, rule_6709, rule_6710, rule_6711, rule_6712, rule_6713, rule_6714, rule_6715, rule_6716, rule_6717, rule_6718, rule_6719, rule_6720, rule_6721, rule_6722, rule_6723, rule_6724, rule_6725, rule_6726, rule_6727, rule_6728, rule_6729, rule_6730, rule_6731, rule_6732, rule_6733, rule_6734, rule_6735, rule_6736, rule_6737, rule_6738, rule_6739, rule_6740, rule_6741, rule_6742, rule_6743, rule_6744, rule_6745, rule_6746, rule_6747, rule_6748, rule_6749, rule_6750, rule_6751, rule_6752, rule_6753, rule_6754, rule_6755, rule_6756, rule_6757, rule_6758, rule_6759, rule_6760, rule_6761, rule_6762, rule_6763, rule_6764, rule_6765, rule_6766, rule_6767, rule_6768, rule_6769, rule_6770, rule_6771, rule_6772, rule_6773, rule_6774, rule_6775, rule_6776, rule_6777, rule_6778, rule_6779, rule_6780, rule_6781, rule_6782, rule_6783, rule_6784, rule_6785, rule_6786, rule_6787, rule_6788, rule_6789, rule_6790, rule_6791, rule_6792, rule_6793, rule_6794, rule_6795, rule_6796, rule_6797, rule_6798, rule_6799, rule_6800, rule_6801, rule_6802, rule_6803, rule_6804, rule_6805, rule_6806, rule_6807, rule_6808, rule_6809, rule_6810, rule_6811, rule_6812, rule_6813, rule_6814, rule_6815, rule_6816, rule_6817, rule_6818, rule_6819, rule_6820, rule_6821, rule_6822, rule_6823, rule_6824, rule_6825, rule_6826, rule_6827, rule_6828, rule_6829, rule_6830, rule_6831, rule_6832, rule_6833, rule_6834, rule_6835, rule_6836, rule_6837, rule_6838, rule_6839, rule_6840, rule_6841, rule_6842, rule_6843, rule_6844, rule_6845, rule_6846, rule_6847, rule_6848, rule_6849, rule_6850, rule_6851, rule_6852, rule_6853, rule_6854, rule_6855, rule_6856, rule_6857, rule_6858, rule_6859, rule_6860, rule_6861, rule_6862, rule_6863, rule_6864, rule_6865, rule_6866, rule_6867, rule_6868, rule_6869, rule_6870, rule_6871, rule_6872, rule_6873, rule_6874, rule_6875, rule_6876, rule_6877, rule_6878, rule_6879, rule_6880, rule_6881, rule_6882, rule_6883, rule_6884, rule_6885, rule_6886, rule_6887, rule_6888, rule_6889, rule_6890, rule_6891, rule_6892, rule_6893, rule_6894, rule_6895, rule_6896, rule_6897, rule_6898, rule_6899, rule_6900, rule_6901, rule_6902, rule_6903, rule_6904, rule_6905, rule_6906, rule_6907, rule_6908, rule_6909, rule_6910, rule_6911, rule_6912, rule_6913, rule_6914, rule_6915, rule_6916, rule_6917, rule_6918, rule_6919, rule_6920, rule_6921, rule_6922, rule_6923, rule_6924, rule_6925, rule_6926, rule_6927, rule_6928, rule_6929, rule_6930, rule_6931, rule_6932, rule_6933, rule_6934, rule_6935, rule_6936, rule_6937, rule_6938, rule_6939, rule_6940, rule_6941, rule_6942, rule_6943, rule_6944, rule_6945, rule_6946, rule_6947, rule_6948, rule_6949, rule_6950, rule_6951, rule_6952, rule_6953, rule_6954, rule_6955, rule_6956, rule_6957, rule_6958, rule_6959, rule_6960, rule_6961, rule_6962, rule_6963, rule_6964, rule_6965, rule_6966, rule_6967, rule_6968, rule_6969, rule_6970, rule_6971, rule_6972, rule_6973, rule_6974, rule_6975, rule_6976, rule_6977, rule_6978, rule_6979, rule_6980, rule_6981, rule_6982, rule_6983, rule_6984, rule_6985, rule_6986, rule_6987, rule_6988, rule_6989, rule_6990, rule_6991, rule_6992, rule_6993, rule_6994, rule_6995, rule_6996, rule_6997, rule_6998, rule_6999, rule_7000, rule_7001, rule_7002, rule_7003, rule_7004, rule_7005, rule_7006, rule_7007, rule_7008, rule_7009, rule_7010, rule_7011, rule_7012, rule_7013, rule_7014, rule_7015, rule_7016, rule_7017, rule_7018, rule_7019, rule_7020, rule_7021, rule_7022, rule_7023, rule_7024, rule_7025, rule_7026, rule_7027, rule_7028, rule_7029, rule_7030, rule_7031, rule_7032, rule_7033, rule_7034, rule_7035, rule_7036, rule_7037, rule_7038, rule_7039, rule_7040, rule_7041, rule_7042, rule_7043, rule_7044, rule_7045, rule_7046, rule_7047, rule_7048, rule_7049, rule_7050, rule_7051, rule_7052, rule_7053, rule_7054, rule_7055, rule_7056, rule_7057, rule_7058, rule_7059, rule_7060, rule_7061, rule_7062, rule_7063, rule_7064, rule_7065, rule_7066, rule_7067, rule_7068, rule_7069, rule_7070, rule_7071, rule_7072, rule_7073, rule_7074, rule_7075, rule_7076, rule_7077, rule_7078, rule_7079, rule_7080, rule_7081, rule_7082, rule_7083, rule_7084, rule_7085, rule_7086, rule_7087, rule_7088, rule_7089, rule_7090, rule_7091, rule_7092, rule_7093, rule_7094, rule_7095, rule_7096, rule_7097, rule_7098, rule_7099, rule_7100, rule_7101, rule_7102, rule_7103, rule_7104, rule_7105, rule_7106, rule_7107, rule_7108, rule_7109, rule_7110, rule_7111, rule_7112, rule_7113, rule_7114, rule_7115, rule_7116, rule_7117, rule_7118, rule_7119, rule_7120, rule_7121, rule_7122, rule_7123, rule_7124, rule_7125, rule_7126, rule_7127, rule_7128, rule_7129, rule_7130, rule_7131, rule_7132, rule_7133, rule_7134, rule_7135, rule_7136, rule_7137, rule_7138, rule_7139, rule_7140, rule_7141, rule_7142, rule_7143, rule_7144, rule_7145, rule_7146, rule_7147, rule_7148, rule_7149, rule_7150, rule_7151, rule_7152, rule_7153, rule_7154, rule_7155, rule_7156, rule_7157, rule_7158, rule_7159, rule_7160, rule_7161, rule_7162, rule_7163, rule_7164, rule_7165, rule_7166, rule_7167, rule_7168, rule_7169, rule_7170, rule_7171, rule_7172, rule_7173, rule_7174, rule_7175, rule_7176, rule_7177, rule_7178, rule_7179, rule_7180, rule_7181, rule_7182, rule_7183, rule_7184, rule_7185, rule_7186, rule_7187, rule_7188, rule_7189, rule_7190, rule_7191, rule_7192, rule_7193, rule_7194, rule_7195, rule_7196, rule_7197, rule_7198, rule_7199, rule_7200, rule_7201, rule_7202, rule_7203, rule_7204, rule_7205, rule_7206, rule_7207, rule_7208, rule_7209, rule_7210, rule_7211, rule_7212, rule_7213, rule_7214, rule_7215, rule_7216, rule_7217, rule_7218, rule_7219, rule_7220, rule_7221, rule_7222, rule_7223, rule_7224, rule_7225, rule_7226, rule_7227, rule_7228, rule_7229, rule_7230, rule_7231, rule_7232, rule_7233, rule_7234, rule_7235, rule_7236, rule_7237, rule_7238, rule_7239, rule_7240, rule_7241, rule_7242, rule_7243, rule_7244, rule_7245, rule_7246, rule_7247, rule_7248, rule_7249, rule_7250, rule_7251, rule_7252, rule_7253, rule_7254, rule_7255, rule_7256, rule_7257, rule_7258, rule_7259, rule_7260, rule_7261, rule_7262, rule_7263, rule_7264, rule_7265, rule_7266, rule_7267, rule_7268, rule_7269, rule_7270, rule_7271, rule_7272, rule_7273, rule_7274, rule_7275, rule_7276, rule_7277, rule_7278, rule_7279, rule_7280, rule_7281, rule_7282, rule_7283, rule_7284, rule_7285, rule_7286, rule_7287, rule_7288, rule_7289, rule_7290, rule_7291, rule_7292, rule_7293, rule_7294, rule_7295, rule_7296, rule_7297, rule_7298, rule_7299, rule_7300, rule_7301, rule_7302, rule_7303, rule_7304, rule_7305, rule_7306, rule_7307, rule_7308, rule_7309, rule_7310, rule_7311, rule_7312, rule_7313, rule_7314, rule_7315, rule_7316, rule_7317, rule_7318, rule_7319, rule_7320, rule_7321, rule_7322, rule_7323, rule_7324, rule_7325, rule_7326, rule_7327, rule_7328, rule_7329, rule_7330, rule_7331, rule_7332, rule_7333, rule_7334, rule_7335, rule_7336, rule_7337, rule_7338, rule_7339, rule_7340, rule_7341, rule_7342, rule_7343, rule_7344, rule_7345, rule_7346, rule_7347, rule_7348, rule_7349, rule_7350, rule_7351, rule_7352, rule_7353, rule_7354, rule_7355, rule_7356, rule_7357, rule_7358, rule_7359, rule_7360, rule_7361, rule_7362, rule_7363, rule_7364, rule_7365, rule_7366, rule_7367, rule_7368, rule_7369, rule_7370, rule_7371, rule_7372, rule_7373, rule_7374, rule_7375, rule_7376, rule_7377, rule_7378, rule_7379, rule_7380, rule_7381, rule_7382, rule_7383, rule_7384, rule_7385, rule_7386, rule_7387, rule_7388, rule_7389, rule_7390, rule_7391, rule_7392, rule_7393, rule_7394, rule_7395, rule_7396, rule_7397, rule_7398, rule_7399, rule_7400, rule_7401, rule_7402, rule_7403, rule_7404, rule_7405, rule_7406, rule_7407, rule_7408, rule_7409, rule_7410, rule_7411, rule_7412, rule_7413, rule_7414, rule_7415, rule_7416, rule_7417, rule_7418, rule_7419, rule_7420, rule_7421, rule_7422, rule_7423, rule_7424, rule_7425, rule_7426, rule_7427, rule_7428, rule_7429, rule_7430, rule_7431, rule_7432, rule_7433, rule_7434, rule_7435, rule_7436, rule_7437, rule_7438, rule_7439, rule_7440, rule_7441, rule_7442, rule_7443, rule_7444, rule_7445, rule_7446, rule_7447, rule_7448, rule_7449, rule_7450, rule_7451, rule_7452, rule_7453, rule_7454, rule_7455, rule_7456, rule_7457, rule_7458, rule_7459, rule_7460, rule_7461, rule_7462, rule_7463, rule_7464, rule_7465, rule_7466, rule_7467, rule_7468, rule_7469, rule_7470, rule_7471, rule_7472, rule_7473, rule_7474, rule_7475, rule_7476, rule_7477, rule_7478, rule_7479, rule_7480, rule_7481, rule_7482, rule_7483, rule_7484, rule_7485, rule_7486, rule_7487, rule_7488, rule_7489, rule_7490, rule_7491, rule_7492, rule_7493, rule_7494, rule_7495, rule_7496, rule_7497, rule_7498, rule_7499, rule_7500, rule_7501, rule_7502, rule_7503, rule_7504, rule_7505, rule_7506, rule_7507, rule_7508, rule_7509, rule_7510, rule_7511, rule_7512, rule_7513, rule_7514, rule_7515, rule_7516, rule_7517, rule_7518, rule_7519, rule_7520, rule_7521, rule_7522, rule_7523, rule_7524, rule_7525, rule_7526, rule_7527, rule_7528, rule_7529, rule_7530, rule_7531, rule_7532, rule_7533, rule_7534, rule_7535, rule_7536, rule_7537, rule_7538, rule_7539, rule_7540, rule_7541, rule_7542, rule_7543, rule_7544, rule_7545, rule_7546, rule_7547, rule_7548, rule_7549, rule_7550, rule_7551, rule_7552, rule_7553, rule_7554, rule_7555, rule_7556, rule_7557, rule_7558, rule_7559, rule_7560, rule_7561, rule_7562, rule_7563, rule_7564, rule_7565, rule_7566, rule_7567, rule_7568, rule_7569, rule_7570, rule_7571, rule_7572, rule_7573, rule_7574, rule_7575, rule_7576, rule_7577, rule_7578, rule_7579, rule_7580, rule_7581, rule_7582, rule_7583, rule_7584, rule_7585, rule_7586, rule_7587, rule_7588, rule_7589, rule_7590, rule_7591, rule_7592, rule_7593, rule_7594, rule_7595, rule_7596, rule_7597, rule_7598, rule_7599, rule_7600, rule_7601, rule_7602, rule_7603, rule_7604, rule_7605, rule_7606, rule_7607, rule_7608, rule_7609, rule_7610, rule_7611, rule_7612, rule_7613, rule_7614, rule_7615, rule_7616, rule_7617, rule_7618, rule_7619, rule_7620, rule_7621, rule_7622, rule_7623, rule_7624, rule_7625, rule_7626, rule_7627, rule_7628, rule_7629, rule_7630, rule_7631, rule_7632, rule_7633, rule_7634, rule_7635, rule_7636, rule_7637, rule_7638, rule_7639, rule_7640, rule_7641, rule_7642, rule_7643, rule_7644, rule_7645, rule_7646, rule_7647, rule_7648, rule_7649, rule_7650, rule_7651, rule_7652, rule_7653, rule_7654, rule_7655, rule_7656, rule_7657, rule_7658, rule_7659, rule_7660, rule_7661, rule_7662, rule_7663, rule_7664, rule_7665, rule_7666, rule_7667, rule_7668, rule_7669, rule_7670, rule_7671, rule_7672, rule_7673, rule_7674, rule_7675, rule_7676, rule_7677, rule_7678, rule_7679, rule_7680, rule_7681, rule_7682, rule_7683, rule_7684, rule_7685, rule_7686, rule_7687, rule_7688, rule_7689, rule_7690, rule_7691, rule_7692, rule_7693, rule_7694, rule_7695, rule_7696, rule_7697, rule_7698, rule_7699, rule_7700, rule_7701, rule_7702, rule_7703, rule_7704, rule_7705, rule_7706, rule_7707, rule_7708, rule_7709, rule_7710, rule_7711, rule_7712, rule_7713, rule_7714, rule_7715, rule_7716, rule_7717, rule_7718, rule_7719, rule_7720, rule_7721, rule_7722, rule_7723, rule_7724, rule_7725, rule_7726, rule_7727, rule_7728, rule_7729, rule_7730, rule_7731, rule_7732, rule_7733, rule_7734, rule_7735, rule_7736, rule_7737, rule_7738, rule_7739, rule_7740, rule_7741, rule_7742, rule_7743, rule_7744, rule_7745, rule_7746, rule_7747, rule_7748, rule_7749, rule_7750, rule_7751, rule_7752, rule_7753, rule_7754, rule_7755, rule_7756, rule_7757, rule_7758, rule_7759, rule_7760, rule_7761, rule_7762, rule_7763, rule_7764, rule_7765, rule_7766, rule_7767, rule_7768, rule_7769, rule_7770, rule_7771, rule_7772, rule_7773, rule_7774, rule_7775, rule_7776, rule_7777, rule_7778, rule_7779, rule_7780, rule_7781, rule_7782, rule_7783, rule_7784, rule_7785, rule_7786, rule_7787, rule_7788, rule_7789, rule_7790, rule_7791, rule_7792, rule_7793, rule_7794, rule_7795, rule_7796, rule_7797, rule_7798, rule_7799, rule_7800, rule_7801, rule_7802, rule_7803, rule_7804, rule_7805, rule_7806, rule_7807, rule_7808, rule_7809, rule_7810, rule_7811, rule_7812, rule_7813, rule_7814, rule_7815, rule_7816, rule_7817, rule_7818, rule_7819, rule_7820, rule_7821, rule_7822, rule_7823, rule_7824, rule_7825, rule_7826, rule_7827, rule_7828, rule_7829, rule_7830, rule_7831, rule_7832, rule_7833, rule_7834, rule_7835, rule_7836, rule_7837, rule_7838, rule_7839, rule_7840, rule_7841, rule_7842, rule_7843, rule_7844, rule_7845, rule_7846, rule_7847, rule_7848, rule_7849, rule_7850, rule_7851, rule_7852, rule_7853, rule_7854, rule_7855, rule_7856, rule_7857, rule_7858, rule_7859, rule_7860, rule_7861, rule_7862, rule_7863, rule_7864, rule_7865, rule_7866, rule_7867, rule_7868, rule_7869, rule_7870, rule_7871, rule_7872, rule_7873, rule_7874, rule_7875, rule_7876, rule_7877, rule_7878, rule_7879, rule_7880, rule_7881, rule_7882, rule_7883, rule_7884, rule_7885, rule_7886, rule_7887, rule_7888, rule_7889, rule_7890, rule_7891, rule_7892, rule_7893, rule_7894, rule_7895, rule_7896, rule_7897, rule_7898, rule_7899, rule_7900, rule_7901, rule_7902, rule_7903, rule_7904, rule_7905, rule_7906, rule_7907, rule_7908, rule_7909, rule_7910, rule_7911, rule_7912, rule_7913, rule_7914, rule_7915, rule_7916, rule_7917, rule_7918, rule_7919, rule_7920, rule_7921, rule_7922, rule_7923, rule_7924, rule_7925, rule_7926, rule_7927, rule_7928, rule_7929, rule_7930, rule_7931, rule_7932, rule_7933, rule_7934, rule_7935, rule_7936, rule_7937, rule_7938, rule_7939, rule_7940, rule_7941, rule_7942, rule_7943, rule_7944, rule_7945, rule_7946, rule_7947, rule_7948, rule_7949, rule_7950, rule_7951, rule_7952" *)
    rule rule_6785;
        ChannelMessage t;
        t <- mod_5532.get(0);
        mod_4633.put(3, t);
    endrule
    rule rule_6786;
        ChannelMessage t;
        t <- mod_5600.get(4);
        mod_164.put(1, t);
    endrule
    rule rule_6787;
        ChannelMessage t;
        t <- mod_5451.get(0);
        mod_1025.put(2, t);
    endrule
    rule rule_6788;
        ChannelMessage t;
        t <- mod_5457.get(0);
        mod_4182.put(4, t);
    endrule
    rule rule_6789;
        ChannelMessage t;
        t <- mod_902.get(0);
        mod_5382.put(0, t);
    endrule
    rule rule_6790;
        ChannelMessage t;
        t <- mod_984.get(0);
        mod_5313.put(103, t);
    endrule
    rule rule_6791;
        ChannelMessage t;
        t <- mod_3321.get(1);
        mod_5313.put(46, t);
    endrule
    rule rule_6792;
        ChannelMessage t;
        t <- mod_5309.get(93);
        mod_3813.put(0, t);
    endrule
    rule rule_6793;
        ChannelMessage t;
        t <- mod_3608.get(3);
        mod_5401.put(0, t);
    endrule
    rule rule_6794;
        ChannelMessage t;
        t <- mod_5565.get(0);
        mod_4633.put(4, t);
    endrule
    rule rule_6795;
        ChannelMessage t;
        t <- mod_5329.get(0);
        mod_1845.put(4, t);
    endrule
    rule rule_6796;
        ChannelMessage t;
        t <- mod_5309.get(55);
        mod_2255.put(0, t);
    endrule
    rule rule_6797;
        ChannelMessage t;
        t <- mod_5402.get(0);
        mod_3690.put(4, t);
    endrule
    rule rule_6798;
        ChannelMessage t;
        t <- mod_5627.get(0);
        mod_4428.put(3, t);
    endrule
    rule rule_6799;
        ChannelMessage t;
        t <- mod_5584.get(0);
        mod_1517.put(3, t);
    endrule
    rule rule_6800;
        ChannelMessage t;
        t <- mod_5648.get(0);
        mod_2460.put(2, t);
    endrule
    rule rule_6801;
        ChannelMessage t;
        t <- mod_5326.get(1);
        mod_5372.put(1, t);
    endrule
    rule rule_6802;
        ChannelMessage t;
        t <- mod_2214.get(3);
        mod_5420.put(0, t);
    endrule
    rule rule_6803;
        ChannelMessage t;
        t <- mod_5309.get(101);
        mod_4141.put(0, t);
    endrule
    rule rule_6804;
        ChannelMessage t;
        t <- mod_1927.get(1);
        mod_5310.put(0, t);
    endrule
    rule rule_6805;
        ChannelMessage t;
        t <- mod_5390.get(0);
        mod_1230.put(4, t);
    endrule
    rule rule_6806;
        ChannelMessage t;
        t <- mod_5364.get(0);
        mod_2255.put(3, t);
    endrule
    rule rule_6807;
        ChannelMessage t;
        t <- mod_5500.get(0);
        mod_123.put(3, t);
    endrule
    rule rule_6808;
        ChannelMessage t;
        t <- mod_5309.get(107);
        mod_4387.put(0, t);
    endrule
    rule rule_6809;
        ChannelMessage t;
        t <- mod_82.get(1);
        mod_5272.put(0, t);
    endrule
    rule rule_6810;
        ChannelMessage t;
        t <- mod_4510.get(3);
        mod_5558.put(0, t);
    endrule
    rule rule_6811;
        ChannelMessage t;
        t <- mod_5600.get(116);
        mod_4756.put(1, t);
    endrule
    rule rule_6812;
        ChannelMessage t;
        t <- mod_1599.get(0);
        mod_5313.put(88, t);
    endrule
    rule rule_6813;
        ChannelMessage t;
        t <- mod_3813.get(1);
        mod_5345.put(0, t);
    endrule
    rule rule_6814;
        ChannelMessage t;
        t <- mod_5496.get(0);
        mod_3731.put(3, t);
    endrule
    rule rule_6815;
        ChannelMessage t;
        t <- mod_5309.get(62);
        mod_2542.put(0, t);
    endrule
    rule rule_6816;
        ChannelMessage t;
        t <- mod_5380.get(0);
        mod_1312.put(3, t);
    endrule
    rule rule_6817;
        ChannelMessage t;
        t <- mod_5461.get(0);
        mod_246.put(3, t);
    endrule
    rule rule_6818;
        ChannelMessage t;
        t <- mod_5309.get(118);
        mod_4838.put(0, t);
    endrule
    rule rule_6819;
        ChannelMessage t;
        t <- mod_5589.get(0);
        mod_1558.put(2, t);
    endrule
    rule rule_6820;
        ChannelMessage t;
        t <- mod_5594.get(0);
        mod_4305.put(4, t);
    endrule
    rule rule_6821;
        ChannelMessage t;
        t <- mod_5309.get(8);
        mod_328.put(0, t);
    endrule
    rule rule_6822;
        ChannelMessage t;
        t <- mod_5408.get(0);
        mod_2952.put(2, t);
    endrule
    rule rule_6823;
        ChannelMessage t;
        t <- mod_5309.get(108);
        mod_4428.put(0, t);
    endrule
    rule rule_6824;
        ChannelMessage t;
        t <- mod_5600.get(64);
        mod_2624.put(1, t);
    endrule
    rule rule_6825;
        ChannelMessage t;
        t <- mod_5600.get(88);
        mod_3608.put(1, t);
    endrule
    rule rule_6826;
        ChannelMessage t;
        t <- mod_5600.get(103);
        mod_4223.put(1, t);
    endrule
    rule rule_6827;
        ChannelMessage t;
        t <- mod_3608.get(0);
        mod_5346.put(0, t);
    endrule
    rule rule_6828;
        ChannelMessage t;
        t <- mod_5600.get(71);
        mod_2911.put(1, t);
    endrule
    rule rule_6829;
        ChannelMessage t;
        t <- mod_5587.get(0);
        mod_1722.put(2, t);
    endrule
    rule rule_6830;
        ChannelMessage t;
        t <- mod_1312.get(3);
        mod_5380.put(0, t);
    endrule
    rule rule_6831;
        ChannelMessage t;
        t <- mod_1353.get(1);
        mod_5471.put(0, t);
    endrule
    rule rule_6832;
        ChannelMessage t;
        t <- mod_5391.get(0);
        mod_4551.put(2, t);
    endrule
    rule rule_6833;
        ChannelMessage t;
        t <- mod_5600.get(87);
        mod_3567.put(1, t);
    endrule
    rule rule_6834;
        ChannelMessage t;
        t <- mod_5309.get(102);
        mod_4182.put(0, t);
    endrule
    rule rule_6835;
        ChannelMessage t;
        t <- mod_861.get(0);
        mod_5313.put(106, t);
    endrule
    rule rule_6836;
        ChannelMessage t;
        t <- mod_2337.get(1);
        mod_5313.put(70, t);
    endrule
    rule rule_6837;
        ChannelMessage t;
        t <- mod_5600.get(36);
        mod_1476.put(1, t);
    endrule
    rule rule_6838;
        ChannelMessage t;
        t <- mod_5646.get(0);
        mod_5166.put(4, t);
    endrule
    rule rule_6839;
        ChannelMessage t;
        t <- mod_5600.get(33);
        mod_1353.put(1, t);
    endrule
    rule rule_6840;
        ChannelMessage t;
        t <- mod_984.get(3);
        mod_5353.put(0, t);
    endrule
    rule rule_6841;
        ChannelMessage t;
        t <- mod_5600.get(28);
        mod_1148.put(1, t);
    endrule
    rule rule_6842;
        ChannelMessage t;
        t <- mod_1435.get(0);
        mod_5417.put(0, t);
    endrule
    rule rule_6843;
        ChannelMessage t;
        t <- mod_5309.get(115);
        mod_4715.put(0, t);
    endrule
    rule rule_6844;
        ChannelMessage t;
        t <- mod_5624.get(0);
        mod_1025.put(3, t);
    endrule
    rule rule_6845;
        ChannelMessage t;
        t <- mod_5600.get(68);
        mod_2788.put(1, t);
    endrule
    rule rule_6846;
        ChannelMessage t;
        t <- mod_4797.get(0);
        mod_5354.put(0, t);
    endrule
    rule rule_6847;
        ChannelMessage t;
        t <- mod_4838.get(0);
        mod_5313.put(9, t);
    endrule
    rule rule_6848;
        ChannelMessage t;
        t <- mod_410.get(3);
        mod_5313.put(117, t);
    endrule
    rule rule_6849;
        ChannelMessage t;
        t <- mod_5465.get(0);
        mod_1230.put(3, t);
    endrule
    rule rule_6850;
        ChannelMessage t;
        t <- mod_5600.get(80);
        mod_3280.put(1, t);
    endrule
    rule rule_6851;
        ChannelMessage t;
        t <- mod_5600.get(37);
        mod_1517.put(1, t);
    endrule
    rule rule_6852;
        ChannelMessage t;
        t <- mod_3280.get(0);
        mod_5313.put(47, t);
    endrule
    rule rule_6853;
        ChannelMessage t;
        t <- mod_3813.get(2);
        mod_5361.put(0, t);
    endrule
    rule rule_6854;
        ChannelMessage t;
        t <- mod_3567.get(0);
        mod_5606.put(0, t);
    endrule
    rule rule_6855;
        ChannelMessage t;
        t <- mod_5288.get(0);
        mod_3895.put(3, t);
    endrule
    rule rule_6856;
        ChannelMessage t;
        t <- mod_5562.get(0);
        mod_4018.put(2, t);
    endrule
    rule rule_6857;
        ChannelMessage t;
        t <- mod_5600.get(48);
        mod_1968.put(1, t);
    endrule
    rule rule_6858;
        ChannelMessage t;
        t <- mod_5426.get(0);
        mod_5523.put(0, t);
    endrule
    rule rule_6859;
        ChannelMessage t;
        t <- mod_5579.get(0);
        mod_1394.put(3, t);
    endrule
    rule rule_6860;
        ChannelMessage t;
        t <- mod_5600.get(8);
        mod_328.put(1, t);
    endrule
    rule rule_6861;
        ChannelMessage t;
        t <- mod_3321.get(0);
        mod_5641.put(0, t);
    endrule
    rule rule_6862;
        ChannelMessage t;
        t <- mod_574.get(3);
        mod_5517.put(0, t);
    endrule
    rule rule_6863;
        ChannelMessage t;
        t <- mod_5600.get(73);
        mod_2993.put(1, t);
    endrule
    rule rule_6864;
        ChannelMessage t;
        t <- mod_5600.get(110);
        mod_4510.put(1, t);
    endrule
    rule rule_6865;
        ChannelMessage t;
        t <- mod_5600.get(50);
        mod_2050.put(1, t);
    endrule
    rule rule_6866;
        ChannelMessage t;
        t <- mod_4346.get(0);
        mod_5439.put(0, t);
    endrule
    rule rule_6867;
        ChannelMessage t;
        t <- mod_5309.get(91);
        mod_3731.put(0, t);
    endrule
    rule rule_6868;
        ChannelMessage t;
        t <- mod_5419.get(0);
        mod_902.put(2, t);
    endrule
    rule rule_6869;
        ChannelMessage t;
        t <- mod_3485.get(3);
        mod_5400.put(0, t);
    endrule
    rule rule_6870;
        ChannelMessage t;
        t <- mod_3813.get(3);
        mod_5313.put(34, t);
    endrule
    rule rule_6871;
        ChannelMessage t;
        t <- mod_5125.get(0);
        mod_5313.put(2, t);
    endrule
    rule rule_6872;
        ChannelMessage t;
        t <- mod_5309.get(22);
        mod_902.put(0, t);
    endrule
    rule rule_6873;
        ChannelMessage t;
        t <- mod_3608.get(2);
        mod_5303.put(0, t);
    endrule
    rule rule_6874;
        ChannelMessage t;
        t <- mod_5309.get(63);
        mod_2583.put(0, t);
    endrule
    rule rule_6875;
        ChannelMessage t;
        t <- mod_5309.get(72);
        mod_2952.put(0, t);
    endrule
    rule rule_6876;
        ChannelMessage t;
        t <- mod_5311.get(0);
        mod_328.put(2, t);
    endrule
    rule rule_6877;
        ChannelMessage t;
        t <- mod_5492.get(0);
        mod_4633.put(2, t);
    endrule
    rule rule_6878;
        ChannelMessage t;
        t <- mod_1722.get(0);
        mod_5611.put(0, t);
    endrule
    rule rule_6879;
        ChannelMessage t;
        t <- mod_5600.get(21);
        mod_861.put(1, t);
    endrule
    rule rule_6880;
        ChannelMessage t;
        t <- mod_5341.get(0);
        mod_205.put(4, t);
    endrule
    rule rule_6881;
        ChannelMessage t;
        t <- mod_5600.get(94);
        mod_3854.put(1, t);
    endrule
    rule rule_6882;
        ChannelMessage t;
        t <- mod_5600.get(118);
        mod_4838.put(1, t);
    endrule
    rule rule_6883;
        ChannelMessage t;
        t <- mod_5608.get(0);
        mod_2829.put(4, t);
    endrule
    rule rule_6884;
        ChannelMessage t;
        t <- mod_5619.get(0);
        mod_1763.put(2, t);
    endrule
    rule rule_6885;
        ChannelMessage t;
        t <- mod_5084.get(2);
        mod_5313.put(3, t);
    endrule
    rule rule_6886;
        ChannelMessage t;
        t <- mod_5610.get(0);
        mod_492.put(4, t);
    endrule
    rule rule_6887;
        ChannelMessage t;
        t <- mod_1312.get(0);
        mod_5313.put(95, t);
    endrule
    rule rule_6888;
        ChannelMessage t;
        t <- mod_5309.get(74);
        mod_3034.put(0, t);
    endrule
    rule rule_6889;
        ChannelMessage t;
        t <- mod_5458.get(0);
        mod_4838.put(3, t);
    endrule
    rule rule_6890;
        ChannelMessage t;
        t <- mod_5166.get(2);
        mod_5313.put(1, t);
    endrule
    rule rule_6891;
        ChannelMessage t;
        t <- mod_3936.get(3);
        mod_5280.put(0, t);
    endrule
    rule rule_6892;
        ChannelMessage t;
        t <- mod_5309.get(25);
        mod_1025.put(0, t);
    endrule
    rule rule_6893;
        ChannelMessage t;
        t <- mod_820.get(2);
        mod_5405.put(0, t);
    endrule
    rule rule_6894;
        ChannelMessage t;
        t <- mod_2419.get(2);
        mod_5605.put(0, t);
    endrule
    rule rule_6895;
        ChannelMessage t;
        t <- mod_4920.get(3);
        mod_5536.put(0, t);
    endrule
    rule rule_6896;
        ChannelMessage t;
        t <- mod_5309.get(21);
        mod_861.put(0, t);
    endrule
    rule rule_6897;
        ChannelMessage t;
        t <- mod_5309.get(31);
        mod_1271.put(0, t);
    endrule
    rule rule_6898;
        ChannelMessage t;
        t <- mod_5571.get(0);
        mod_2132.put(4, t);
    endrule
    rule rule_6899;
        ChannelMessage t;
        t <- mod_5490.get(0);
        mod_943.put(4, t);
    endrule
    rule rule_6900;
        ChannelMessage t;
        t <- mod_2296.get(3);
        mod_5270.put(0, t);
    endrule
    rule rule_6901;
        ChannelMessage t;
        t <- mod_3239.get(2);
        mod_5498.put(0, t);
    endrule
    rule rule_6902;
        ChannelMessage t;
        t <- mod_5043.get(0);
        mod_5274.put(0, t);
    endrule
    rule rule_6903;
        ChannelMessage t;
        t <- mod_5600.get(29);
        mod_1189.put(1, t);
    endrule
    rule rule_6904;
        ChannelMessage t;
        t <- mod_4346.get(1);
        mod_5264.put(0, t);
    endrule
    rule rule_6905;
        ChannelMessage t;
        t <- mod_4182.get(1);
        mod_5457.put(0, t);
    endrule
    rule rule_6906;
        ChannelMessage t;
        t <- mod_5309.get(37);
        mod_1517.put(0, t);
    endrule
    rule rule_6907;
        ChannelMessage t;
        t <- mod_5298.get(0);
        mod_697.put(2, t);
    endrule
    rule rule_6908;
        ChannelMessage t;
        t <- mod_4018.get(1);
        mod_5562.put(0, t);
    endrule
    rule rule_6909;
        ChannelMessage t;
        t <- mod_5600.get(86);
        mod_3526.put(1, t);
    endrule
    rule rule_6910;
        ChannelMessage t;
        t <- mod_5309.get(75);
        mod_3075.put(0, t);
    endrule
    rule rule_6911;
        ChannelMessage t;
        t <- mod_4428.get(1);
        mod_5313.put(19, t);
    endrule
    rule rule_6912;
        ChannelMessage t;
        t <- mod_5600.get(60);
        mod_2460.put(1, t);
    endrule
    rule rule_6913;
        ChannelMessage t;
        t <- mod_5414.get(0);
        mod_1476.put(2, t);
    endrule
    rule rule_6914;
        ChannelMessage t;
        t <- mod_5527.get(0);
        mod_1640.put(4, t);
    endrule
    rule rule_6915;
        ChannelMessage t;
        t <- mod_697.get(2);
        mod_5483.put(0, t);
    endrule
    rule rule_6916;
        ChannelMessage t;
        t <- mod_4100.get(1);
        mod_5313.put(27, t);
    endrule
    rule rule_6917;
        ChannelMessage t;
        t <- mod_5600.get(102);
        mod_4182.put(1, t);
    endrule
    rule rule_6918;
        ChannelMessage t;
        t <- mod_5410.get(0);
        mod_4141.put(2, t);
    endrule
    rule rule_6919;
        ChannelMessage t;
        t <- mod_5604.get(0);
        mod_410.put(2, t);
    endrule
    rule rule_6920;
        ChannelMessage t;
        t <- mod_5352.get(0);
        mod_4100.put(2, t);
    endrule
    rule rule_6921;
        ChannelMessage t;
        t <- mod_5309.get(103);
        mod_4223.put(0, t);
    endrule
    rule rule_6922;
        ChannelMessage t;
        t <- mod_5425.get(0);
        mod_4141.put(4, t);
    endrule
    rule rule_6923;
        ChannelMessage t;
        t <- mod_1927.get(2);
        mod_5313.put(80, t);
    endrule
    rule rule_6924;
        ChannelMessage t;
        t <- mod_5600.get(3);
        mod_123.put(1, t);
    endrule
    rule rule_6925;
        ChannelMessage t;
        t <- mod_3772.get(1);
        mod_5313.put(35, t);
    endrule
    rule rule_6926;
        ChannelMessage t;
        t <- mod_5207.get(3);
        mod_5475.put(0, t);
    endrule
    rule rule_6927;
        ChannelMessage t;
        t <- mod_5375.get(0);
        mod_4674.put(2, t);
    endrule
    rule rule_6928;
        ChannelMessage t;
        t <- mod_5600.get(121);
        mod_4961.put(1, t);
    endrule
    rule rule_6929;
        ChannelMessage t;
        t <- mod_5498.get(0);
        mod_3239.put(4, t);
    endrule
    rule rule_6930;
        ChannelMessage t;
        t <- mod_5355.get(0);
        mod_3157.put(4, t);
    endrule
    rule rule_6931;
        ChannelMessage t;
        t <- mod_328.get(3);
        mod_5313.put(119, t);
    endrule
    rule rule_6932;
        ChannelMessage t;
        t <- mod_1107.get(1);
        mod_5299.put(0, t);
    endrule
    rule rule_6933;
        ChannelMessage t;
        t <- mod_5545.get(0);
        mod_2050.put(2, t);
    endrule
    rule rule_6934;
        ChannelMessage t;
        t <- mod_5309.get(29);
        mod_1189.put(0, t);
    endrule
    rule rule_6935;
        ChannelMessage t;
        t <- mod_2501.get(0);
        mod_5369.put(0, t);
    endrule
    rule rule_6936;
        ChannelMessage t;
        t <- mod_3075.get(2);
        mod_5585.put(0, t);
    endrule
    rule rule_6937;
        ChannelMessage t;
        t <- mod_5309.get(11);
        mod_451.put(0, t);
    endrule
    rule rule_6938;
        ChannelMessage t;
        t <- mod_5600.get(22);
        mod_902.put(1, t);
    endrule
    rule rule_6939;
        ChannelMessage t;
        t <- mod_5600.get(59);
        mod_2419.put(1, t);
    endrule
    rule rule_6940;
        ChannelMessage t;
        t <- mod_5455.get(0);
        mod_574.put(3, t);
    endrule
    rule rule_6941;
        ChannelMessage t;
        t <- mod_5596.get(0);
        mod_3403.put(2, t);
    endrule
    rule rule_6942;
        ChannelMessage t;
        t <- mod_1517.get(0);
        mod_5535.put(0, t);
    endrule
    rule rule_6943;
        ChannelMessage t;
        t <- mod_574.get(0);
        mod_5385.put(0, t);
    endrule
    rule rule_6944;
        ChannelMessage t;
        t <- mod_2050.get(3);
        mod_5545.put(0, t);
    endrule
    rule rule_6945;
        ChannelMessage t;
        t <- mod_4346.get(2);
        mod_5520.put(0, t);
    endrule
    rule rule_6946;
        ChannelMessage t;
        t <- mod_1271.get(0);
        mod_5386.put(0, t);
    endrule
    rule rule_6947;
        ChannelMessage t;
        t <- mod_3034.get(3);
        mod_5636.put(0, t);
    endrule
    rule rule_6948;
        ChannelMessage t;
        t <- mod_5309.get(121);
        mod_4961.put(0, t);
    endrule
    rule rule_6949;
        ChannelMessage t;
        t <- mod_3239.get(0);
        mod_5313.put(48, t);
    endrule
    rule rule_6950;
        ChannelMessage t;
        t <- mod_4797.get(3);
        mod_5638.put(0, t);
    endrule
    rule rule_6951;
        ChannelMessage t;
        t <- mod_1148.get(1);
        mod_5313.put(99, t);
    endrule
    rule rule_6952;
        ChannelMessage t;
        t <- mod_5394.get(0);
        mod_287.put(4, t);
    endrule
    rule rule_6953;
        ChannelMessage t;
        t <- mod_5469.get(0);
        mod_2747.put(3, t);
    endrule
    rule rule_6954;
        ChannelMessage t;
        t <- mod_4797.get(2);
        mod_5313.put(10, t);
    endrule
    rule rule_6955;
        ChannelMessage t;
        t <- mod_82.get(3);
        mod_5555.put(0, t);
    endrule
    rule rule_6956;
        ChannelMessage t;
        t <- mod_5580.get(0);
        mod_5309.put(0, t);
    endrule
    rule rule_6957;
        ChannelMessage t;
        t <- mod_2255.get(3);
        mod_5563.put(0, t);
    endrule
    rule rule_6958;
        ChannelMessage t;
        t <- mod_5254.get(0);
        mod_287.put(3, t);
    endrule
    rule rule_6959;
        ChannelMessage t;
        t <- mod_5166.get(1);
        mod_5640.put(0, t);
    endrule
    rule rule_6960;
        ChannelMessage t;
        t <- mod_5516.get(0);
        mod_2583.put(4, t);
    endrule
    rule rule_6961;
        ChannelMessage t;
        t <- mod_5600.get(34);
        mod_1394.put(1, t);
    endrule
    rule rule_6962;
        ChannelMessage t;
        t <- mod_4305.get(2);
        mod_5313.put(22, t);
    endrule
    rule rule_6963;
        ChannelMessage t;
        t <- mod_5378.get(0);
        mod_2952.put(3, t);
    endrule
    rule rule_6964;
        ChannelMessage t;
        t <- mod_5600.get(83);
        mod_3403.put(1, t);
    endrule
    rule rule_6965;
        ChannelMessage t;
        t <- mod_4756.get(2);
        mod_5313.put(11, t);
    endrule
    rule rule_6966;
        ChannelMessage t;
        t <- mod_5459.get(0);
        mod_4223.put(2, t);
    endrule
    rule rule_6967;
        ChannelMessage t;
        t <- mod_1599.get(1);
        mod_5578.put(0, t);
    endrule
    rule rule_6968;
        ChannelMessage t;
        t <- mod_779.get(2);
        mod_5484.put(0, t);
    endrule
    rule rule_6969;
        ChannelMessage t;
        t <- mod_5309.get(12);
        mod_492.put(0, t);
    endrule
    rule rule_6970;
        ChannelMessage t;
        t <- mod_738.get(1);
        mod_5307.put(0, t);
    endrule
    rule rule_6971;
        ChannelMessage t;
        t <- mod_5543.get(0);
        mod_3116.put(2, t);
    endrule
    rule rule_6972;
        ChannelMessage t;
        t <- mod_5463.get(0);
        mod_3526.put(2, t);
    endrule
    rule rule_6973;
        ChannelMessage t;
        t <- mod_4387.get(0);
        mod_5263.put(0, t);
    endrule
    rule rule_6974;
        ChannelMessage t;
        t <- mod_5600.get(74);
        mod_3034.put(1, t);
    endrule
    rule rule_6975;
        ChannelMessage t;
        t <- mod_5314.get(0);
        mod_1517.put(4, t);
    endrule
    rule rule_6976;
        ChannelMessage t;
        t <- mod_5318.get(0);
        mod_2173.put(4, t);
    endrule
    rule rule_6977;
        ChannelMessage t;
        t <- mod_4592.get(2);
        mod_5539.put(0, t);
    endrule
    rule rule_6978;
        ChannelMessage t;
        t <- mod_5302.get(0);
        mod_3362.put(4, t);
    endrule
    rule rule_6979;
        ChannelMessage t;
        t <- mod_1968.get(1);
        mod_5582.put(0, t);
    endrule
    rule rule_6980;
        ChannelMessage t;
        t <- mod_4961.get(1);
        mod_5357.put(0, t);
    endrule
    rule rule_6981;
        ChannelMessage t;
        t <- mod_5332.get(0);
        mod_1107.put(3, t);
    endrule
    rule rule_6982;
        ChannelMessage t;
        t <- mod_5338.get(0);
        mod_2460.put(4, t);
    endrule
    rule rule_6983;
        ChannelMessage t;
        t <- mod_5252.get(0);
        mod_3034.put(3, t);
    endrule
    rule rule_6984;
        ChannelMessage t;
        t <- mod_2706.get(1);
        mod_5268.put(0, t);
    endrule
    rule rule_6985;
        ChannelMessage t;
        t <- mod_5626.get(0);
        mod_5207.put(4, t);
    endrule
    rule rule_6986;
        ChannelMessage t;
        t <- mod_1230.get(1);
        mod_5465.put(0, t);
    endrule
    rule rule_6987;
        ChannelMessage t;
        t <- mod_902.get(1);
        mod_5313.put(105, t);
    endrule
    rule rule_6988;
        ChannelMessage t;
        t <- mod_492.get(1);
        mod_5477.put(0, t);
    endrule
    rule rule_6989;
        ChannelMessage t;
        t <- mod_5510.get(0);
        mod_2173.put(2, t);
    endrule
    rule rule_6990;
        ChannelMessage t;
        t <- mod_5600.get(0);
        mod_0.put(1, t);
    endrule
    rule rule_6991;
        ChannelMessage t;
        t <- mod_164.get(2);
        mod_5566.put(0, t);
    endrule
    rule rule_6992;
        ChannelMessage t;
        t <- mod_5600.get(40);
        mod_1640.put(1, t);
    endrule
    rule rule_6993;
        ChannelMessage t;
        t <- mod_1845.get(2);
        mod_5411.put(0, t);
    endrule
    rule rule_6994;
        ChannelMessage t;
        t <- mod_3116.get(1);
        mod_5470.put(0, t);
    endrule
    rule rule_6995;
        ChannelMessage t;
        t <- mod_2419.get(0);
        mod_5537.put(0, t);
    endrule
    rule rule_6996;
        ChannelMessage t;
        t <- mod_5309.get(27);
        mod_1107.put(0, t);
    endrule
    rule rule_6997;
        ChannelMessage t;
        t <- mod_3403.get(1);
        mod_5313.put(44, t);
    endrule
    rule rule_6998;
        ChannelMessage t;
        t <- mod_5370.get(0);
        mod_656.put(3, t);
    endrule
    rule rule_6999;
        ChannelMessage t;
        t <- mod_5002.get(0);
        mod_5313.put(5, t);
    endrule
    rule rule_7000;
        ChannelMessage t;
        t <- mod_5599.get(0);
        mod_369.put(4, t);
    endrule
    rule rule_7001;
        ChannelMessage t;
        t <- mod_2829.get(3);
        mod_5287.put(0, t);
    endrule
    rule rule_7002;
        ChannelMessage t;
        t <- mod_4264.get(2);
        mod_5389.put(0, t);
    endrule
    rule rule_7003;
        ChannelMessage t;
        t <- mod_4428.get(3);
        mod_5633.put(0, t);
    endrule
    rule rule_7004;
        ChannelMessage t;
        t <- mod_451.get(3);
        mod_5473.put(0, t);
    endrule
    rule rule_7005;
        ChannelMessage t;
        t <- mod_5600.get(27);
        mod_1107.put(1, t);
    endrule
    rule rule_7006;
        ChannelMessage t;
        t <- mod_5600.get(56);
        mod_2296.put(1, t);
    endrule
    rule rule_7007;
        ChannelMessage t;
        t <- mod_984.get(1);
        mod_5335.put(0, t);
    endrule
    rule rule_7008;
        ChannelMessage t;
        t <- mod_5591.get(0);
        mod_2829.put(3, t);
    endrule
    rule rule_7009;
        ChannelMessage t;
        t <- mod_5522.get(0);
        mod_2337.put(3, t);
    endrule
    rule rule_7010;
        ChannelMessage t;
        t <- mod_3526.get(1);
        mod_5463.put(0, t);
    endrule
    rule rule_7011;
        ChannelMessage t;
        t <- mod_4223.get(0);
        mod_5459.put(0, t);
    endrule
    rule rule_7012;
        ChannelMessage t;
        t <- mod_5309.get(32);
        mod_1312.put(0, t);
    endrule
    rule rule_7013;
        ChannelMessage t;
        t <- mod_5309.get(35);
        mod_1435.put(0, t);
    endrule
    rule rule_7014;
        ChannelMessage t;
        t <- mod_5371.get(0);
        mod_2296.put(2, t);
    endrule
    rule rule_7015;
        ChannelMessage t;
        t <- mod_5428.get(0);
        mod_779.put(2, t);
    endrule
    rule rule_7016;
        ChannelMessage t;
        t <- mod_5593.get(0);
        mod_3854.put(2, t);
    endrule
    rule rule_7017;
        ChannelMessage t;
        t <- mod_5278.get(0);
        mod_4756.put(2, t);
    endrule
    rule rule_7018;
        ChannelMessage t;
        t <- mod_5576.get(0);
        mod_3321.put(2, t);
    endrule
    rule rule_7019;
        ChannelMessage t;
        t <- mod_5309.get(4);
        mod_164.put(0, t);
    endrule
    rule rule_7020;
        ChannelMessage t;
        t <- mod_5600.get(108);
        mod_4428.put(1, t);
    endrule
    rule rule_7021;
        ChannelMessage t;
        t <- mod_287.get(3);
        mod_5254.put(0, t);
    endrule
    rule rule_7022;
        ChannelMessage t;
        t <- mod_2747.get(0);
        mod_5313.put(60, t);
    endrule
    rule rule_7023;
        ChannelMessage t;
        t <- mod_5528.get(0);
        mod_0.put(4, t);
    endrule
    rule rule_7024;
        ChannelMessage t;
        t <- mod_5555.get(0);
        mod_82.put(4, t);
    endrule
    rule rule_7025;
        ChannelMessage t;
        t <- mod_5396.get(0);
        mod_4797.put(3, t);
    endrule
    rule rule_7026;
        ChannelMessage t;
        t <- mod_4100.get(3);
        mod_5352.put(0, t);
    endrule
    rule rule_7027;
        ChannelMessage t;
        t <- mod_5600.get(13);
        mod_533.put(1, t);
    endrule
    rule rule_7028;
        ChannelMessage t;
        t <- mod_246.get(3);
        mod_5461.put(0, t);
    endrule
    rule rule_7029;
        ChannelMessage t;
        t <- mod_3444.get(3);
        mod_5494.put(0, t);
    endrule
    rule rule_7030;
        ChannelMessage t;
        t <- mod_2378.get(1);
        mod_5462.put(0, t);
    endrule
    rule rule_7031;
        ChannelMessage t;
        t <- mod_3854.get(2);
        mod_5322.put(0, t);
    endrule
    rule rule_7032;
        ChannelMessage t;
        t <- mod_3362.get(2);
        mod_5313.put(45, t);
    endrule
    rule rule_7033;
        ChannelMessage t;
        t <- mod_5281.get(0);
        mod_3321.put(3, t);
    endrule
    rule rule_7034;
        ChannelMessage t;
        t <- mod_492.get(2);
        mod_5404.put(0, t);
    endrule
    rule rule_7035;
        ChannelMessage t;
        t <- mod_5644.get(0);
        mod_1148.put(2, t);
    endrule
    rule rule_7036;
        ChannelMessage t;
        t <- mod_5282.get(0);
        mod_1640.put(3, t);
    endrule
    rule rule_7037;
        ChannelMessage t;
        t <- mod_3690.get(3);
        mod_5292.put(0, t);
    endrule
    rule rule_7038;
        ChannelMessage t;
        t <- mod_4469.get(0);
        mod_5300.put(0, t);
    endrule
    rule rule_7039;
        ChannelMessage t;
        t <- mod_3239.get(1);
        mod_5534.put(0, t);
    endrule
    rule rule_7040;
        ChannelMessage t;
        t <- mod_3649.get(0);
        mod_5501.put(0, t);
    endrule
    rule rule_7041;
        ChannelMessage t;
        t <- mod_5207.get(2);
        mod_5626.put(0, t);
    endrule
    rule rule_7042;
        ChannelMessage t;
        t <- mod_1599.get(2);
        mod_5257.put(0, t);
    endrule
    rule rule_7043;
        ChannelMessage t;
        t <- mod_5309.get(36);
        mod_1476.put(0, t);
    endrule
    rule rule_7044;
        ChannelMessage t;
        t <- mod_5513.get(0);
        mod_1353.put(2, t);
    endrule
    rule rule_7045;
        ChannelMessage t;
        t <- mod_5600.get(11);
        mod_451.put(1, t);
    endrule
    rule rule_7046;
        ChannelMessage t;
        t <- mod_5477.get(0);
        mod_492.put(3, t);
    endrule
    rule rule_7047;
        ChannelMessage t;
        t <- mod_5600.get(31);
        mod_1271.put(1, t);
    endrule
    rule rule_7048;
        ChannelMessage t;
        t <- mod_2173.get(2);
        mod_5318.put(0, t);
    endrule
    rule rule_7049;
        ChannelMessage t;
        t <- mod_3854.get(0);
        mod_5506.put(0, t);
    endrule
    rule rule_7050;
        ChannelMessage t;
        t <- mod_328.get(2);
        mod_5311.put(0, t);
    endrule
    rule rule_7051;
        ChannelMessage t;
        t <- mod_4182.get(3);
        mod_5609.put(0, t);
    endrule
    rule rule_7052;
        ChannelMessage t;
        t <- mod_5125.get(1);
        mod_5632.put(0, t);
    endrule
    rule rule_7053;
        ChannelMessage t;
        t <- mod_5358.get(0);
        mod_123.put(4, t);
    endrule
    rule rule_7054;
        ChannelMessage t;
        t <- mod_861.get(2);
        mod_5433.put(0, t);
    endrule
    rule rule_7055;
        ChannelMessage t;
        t <- mod_5309.get(85);
        mod_3485.put(0, t);
    endrule
    rule rule_7056;
        ChannelMessage t;
        t <- mod_5331.get(0);
        mod_1271.put(2, t);
    endrule
    rule rule_7057;
        ChannelMessage t;
        t <- mod_5393.get(0);
        mod_1312.put(4, t);
    endrule
    rule rule_7058;
        ChannelMessage t;
        t <- mod_5600.get(114);
        mod_4674.put(1, t);
    endrule
    rule rule_7059;
        ChannelMessage t;
        t <- mod_1804.get(0);
        mod_5277.put(0, t);
    endrule
    rule rule_7060;
        ChannelMessage t;
        t <- mod_1927.get(0);
        mod_5305.put(0, t);
    endrule
    rule rule_7061;
        ChannelMessage t;
        t <- mod_4592.get(1);
        mod_5427.put(0, t);
    endrule
    rule rule_7062;
        ChannelMessage t;
        t <- mod_5276.get(0);
        mod_4920.put(4, t);
    endrule
    rule rule_7063;
        ChannelMessage t;
        t <- mod_5309.get(120);
        mod_4920.put(0, t);
    endrule
    rule rule_7064;
        ChannelMessage t;
        t <- mod_5600.get(123);
        mod_5043.put(1, t);
    endrule
    rule rule_7065;
        ChannelMessage t;
        t <- mod_1476.get(2);
        mod_5581.put(0, t);
    endrule
    rule rule_7066;
        ChannelMessage t;
        t <- mod_4756.get(3);
        mod_5616.put(0, t);
    endrule
    rule rule_7067;
        ChannelMessage t;
        t <- mod_5309.get(20);
        mod_820.put(0, t);
    endrule
    rule rule_7068;
        ChannelMessage t;
        t <- mod_5309.get(98);
        mod_4018.put(0, t);
    endrule
    rule rule_7069;
        ChannelMessage t;
        t <- mod_5600.get(96);
        mod_3936.put(1, t);
    endrule
    rule rule_7070;
        ChannelMessage t;
        t <- mod_5309.get(94);
        mod_3854.put(0, t);
    endrule
    rule rule_7071;
        ChannelMessage t;
        t <- mod_5586.get(0);
        mod_3280.put(4, t);
    endrule
    rule rule_7072;
        ChannelMessage t;
        t <- mod_369.get(0);
        mod_5424.put(0, t);
    endrule
    rule rule_7073;
        ChannelMessage t;
        t <- mod_5600.get(76);
        mod_3116.put(1, t);
    endrule
    rule rule_7074;
        ChannelMessage t;
        t <- mod_5600.get(112);
        mod_4592.put(1, t);
    endrule
    rule rule_7075;
        ChannelMessage t;
        t <- mod_3280.get(1);
        mod_5295.put(0, t);
    endrule
    rule rule_7076;
        ChannelMessage t;
        t <- mod_5296.get(0);
        mod_984.put(4, t);
    endrule
    rule rule_7077;
        ChannelMessage t;
        t <- mod_2788.get(1);
        mod_5313.put(59, t);
    endrule
    rule rule_7078;
        ChannelMessage t;
        t <- mod_5600.get(82);
        mod_3362.put(1, t);
    endrule
    rule rule_7079;
        ChannelMessage t;
        t <- mod_5309.get(64);
        mod_2624.put(0, t);
    endrule
    rule rule_7080;
        ChannelMessage t;
        t <- mod_2009.get(2);
        mod_5313.put(78, t);
    endrule
    rule rule_7081;
        ChannelMessage t;
        t <- mod_3977.get(0);
        mod_5625.put(0, t);
    endrule
    rule rule_7082;
        ChannelMessage t;
        t <- mod_5512.get(0);
        mod_4387.put(2, t);
    endrule
    rule rule_7083;
        ChannelMessage t;
        t <- mod_615.get(0);
        mod_5343.put(0, t);
    endrule
    rule rule_7084;
        ChannelMessage t;
        t <- mod_5345.get(0);
        mod_3813.put(4, t);
    endrule
    rule rule_7085;
        ChannelMessage t;
        t <- mod_4961.get(2);
        mod_5313.put(6, t);
    endrule
    rule rule_7086;
        ChannelMessage t;
        t <- mod_5291.get(0);
        mod_2132.put(2, t);
    endrule
    rule rule_7087;
        ChannelMessage t;
        t <- mod_2501.get(2);
        mod_5541.put(0, t);
    endrule
    rule rule_7088;
        ChannelMessage t;
        t <- mod_2911.get(3);
        mod_5518.put(0, t);
    endrule
    rule rule_7089;
        ChannelMessage t;
        t <- mod_1640.get(2);
        mod_5527.put(0, t);
    endrule
    rule rule_7090;
        ChannelMessage t;
        t <- mod_1230.get(3);
        mod_5313.put(97, t);
    endrule
    rule rule_7091;
        ChannelMessage t;
        t <- mod_5273.get(0);
        mod_2788.put(4, t);
    endrule
    rule rule_7092;
        ChannelMessage t;
        t <- mod_5600.get(44);
        mod_1804.put(1, t);
    endrule
    rule rule_7093;
        ChannelMessage t;
        t <- mod_1886.get(2);
        mod_5313.put(81, t);
    endrule
    rule rule_7094;
        ChannelMessage t;
        t <- mod_5415.get(0);
        mod_2993.put(3, t);
    endrule
    rule rule_7095;
        ChannelMessage t;
        t <- mod_5529.get(0);
        mod_5084.put(3, t);
    endrule
    rule rule_7096;
        ChannelMessage t;
        t <- mod_3895.get(1);
        mod_5313.put(32, t);
    endrule
    rule rule_7097;
        ChannelMessage t;
        t <- mod_5334.get(0);
        mod_943.put(2, t);
    endrule
    rule rule_7098;
        ChannelMessage t;
        t <- mod_5294.get(0);
        mod_4920.put(2, t);
    endrule
    rule rule_7099;
        ChannelMessage t;
        t <- mod_3198.get(1);
        mod_5383.put(0, t);
    endrule
    rule rule_7100;
        ChannelMessage t;
        t <- mod_5320.get(0);
        mod_4674.put(4, t);
    endrule
    rule rule_7101;
        ChannelMessage t;
        t <- mod_5309.get(105);
        mod_4305.put(0, t);
    endrule
    rule rule_7102;
        ChannelMessage t;
        t <- mod_5292.get(0);
        mod_3690.put(3, t);
    endrule
    rule rule_7103;
        ChannelMessage t;
        t <- mod_1681.get(0);
        mod_5568.put(0, t);
    endrule
    rule rule_7104;
        ChannelMessage t;
        t <- mod_1107.get(2);
        mod_5434.put(0, t);
    endrule
    rule rule_7105;
        ChannelMessage t;
        t <- mod_656.get(0);
        mod_5313.put(111, t);
    endrule
    rule rule_7106;
        ChannelMessage t;
        t <- mod_3977.get(1);
        mod_5313.put(30, t);
    endrule
    rule rule_7107;
        ChannelMessage t;
        t <- mod_3444.get(1);
        mod_5313.put(43, t);
    endrule
    rule rule_7108;
        ChannelMessage t;
        t <- mod_5637.get(0);
        mod_3034.put(2, t);
    endrule
    rule rule_7109;
        ChannelMessage t;
        t <- mod_246.get(1);
        mod_5313.put(121, t);
    endrule
    rule rule_7110;
        ChannelMessage t;
        t <- mod_5600.get(125);
        mod_5125.put(1, t);
    endrule
    rule rule_7111;
        ChannelMessage t;
        t <- mod_5487.get(0);
        mod_3731.put(4, t);
    endrule
    rule rule_7112;
        ChannelMessage t;
        t <- mod_5600.get(84);
        mod_3444.put(1, t);
    endrule
    rule rule_7113;
        ChannelMessage t;
        t <- mod_5309.get(7);
        mod_287.put(0, t);
    endrule
    rule rule_7114;
        ChannelMessage t;
        t <- mod_3280.get(3);
        mod_5556.put(0, t);
    endrule
    rule rule_7115;
        ChannelMessage t;
        t <- mod_2132.get(2);
        mod_5533.put(0, t);
    endrule
    rule rule_7116;
        ChannelMessage t;
        t <- mod_205.get(3);
        mod_5359.put(0, t);
    endrule
    rule rule_7117;
        ChannelMessage t;
        t <- mod_451.get(1);
        mod_5480.put(0, t);
    endrule
    rule rule_7118;
        ChannelMessage t;
        t <- mod_3485.get(1);
        mod_5618.put(0, t);
    endrule
    rule rule_7119;
        ChannelMessage t;
        t <- mod_984.get(2);
        mod_5296.put(0, t);
    endrule
    rule rule_7120;
        ChannelMessage t;
        t <- mod_2870.get(2);
        mod_5435.put(0, t);
    endrule
    rule rule_7121;
        ChannelMessage t;
        t <- mod_5600.get(95);
        mod_3895.put(1, t);
    endrule
    rule rule_7122;
        ChannelMessage t;
        t <- mod_2624.get(2);
        mod_5615.put(0, t);
    endrule
    rule rule_7123;
        ChannelMessage t;
        t <- mod_5641.get(0);
        mod_3321.put(4, t);
    endrule
    rule rule_7124;
        ChannelMessage t;
        t <- mod_369.get(3);
        mod_5313.put(118, t);
    endrule
    rule rule_7125;
        ChannelMessage t;
        t <- mod_5309.get(10);
        mod_410.put(0, t);
    endrule
    rule rule_7126;
        ChannelMessage t;
        t <- mod_4592.get(0);
        mod_5313.put(15, t);
    endrule
    rule rule_7127;
        ChannelMessage t;
        t <- mod_4879.get(2);
        mod_5313.put(8, t);
    endrule
    rule rule_7128;
        ChannelMessage t;
        t <- mod_5043.get(1);
        mod_5486.put(0, t);
    endrule
    rule rule_7129;
        ChannelMessage t;
        t <- mod_5309.get(43);
        mod_1763.put(0, t);
    endrule
    rule rule_7130;
        ChannelMessage t;
        t <- mod_533.get(3);
        mod_5313.put(114, t);
    endrule
    rule rule_7131;
        ChannelMessage t;
        t <- mod_697.get(3);
        mod_5313.put(110, t);
    endrule
    rule rule_7132;
        ChannelMessage t;
        t <- mod_5600.get(46);
        mod_1886.put(1, t);
    endrule
    rule rule_7133;
        ChannelMessage t;
        t <- mod_5308.get(0);
        mod_1066.put(4, t);
    endrule
    rule rule_7134;
        ChannelMessage t;
        t <- mod_5601.get(0);
        mod_656.put(2, t);
    endrule
    rule rule_7135;
        ChannelMessage t;
        t <- mod_5605.get(0);
        mod_2419.put(4, t);
    endrule
    rule rule_7136;
        ChannelMessage t;
        t <- mod_4223.get(3);
        mod_5643.put(0, t);
    endrule
    rule rule_7137;
        ChannelMessage t;
        t <- mod_4961.get(3);
        mod_5505.put(0, t);
    endrule
    rule rule_7138;
        ChannelMessage t;
        t <- mod_5600.get(78);
        mod_3198.put(1, t);
    endrule
    rule rule_7139;
        ChannelMessage t;
        t <- mod_5600.get(66);
        mod_2706.put(1, t);
    endrule
    rule rule_7140;
        ChannelMessage t;
        t <- mod_5303.get(0);
        mod_3608.put(3, t);
    endrule
    rule rule_7141;
        ChannelMessage t;
        t <- mod_5600.get(92);
        mod_3772.put(1, t);
    endrule
    rule rule_7142;
        ChannelMessage t;
        t <- mod_5424.get(0);
        mod_369.put(2, t);
    endrule
    rule rule_7143;
        ChannelMessage t;
        t <- mod_5454.get(0);
        mod_2870.put(3, t);
    endrule
    rule rule_7144;
        ChannelMessage t;
        t <- mod_1435.get(1);
        mod_5367.put(0, t);
    endrule
    rule rule_7145;
        ChannelMessage t;
        t <- mod_2419.get(1);
        mod_5444.put(0, t);
    endrule
    rule rule_7146;
        ChannelMessage t;
        t <- mod_2993.get(3);
        mod_5412.put(0, t);
    endrule
    rule rule_7147;
        ChannelMessage t;
        t <- mod_3526.get(3);
        mod_5603.put(0, t);
    endrule
    rule rule_7148;
        ChannelMessage t;
        t <- mod_3567.get(3);
        mod_5315.put(0, t);
    endrule
    rule rule_7149;
        ChannelMessage t;
        t <- mod_5505.get(0);
        mod_4961.put(4, t);
    endrule
    rule rule_7150;
        ChannelMessage t;
        t <- mod_5309.get(59);
        mod_2419.put(0, t);
    endrule
    rule rule_7151;
        ChannelMessage t;
        t <- mod_3772.get(3);
        mod_5612.put(0, t);
    endrule
    rule rule_7152;
        ChannelMessage t;
        t <- mod_1968.get(0);
        mod_5313.put(79, t);
    endrule
    rule rule_7153;
        ChannelMessage t;
        t <- mod_5309.get(28);
        mod_1148.put(0, t);
    endrule
    rule rule_7154;
        ChannelMessage t;
        t <- mod_820.get(1);
        mod_5339.put(0, t);
    endrule
    rule rule_7155;
        ChannelMessage t;
        t <- mod_5600.get(6);
        mod_246.put(1, t);
    endrule
    rule rule_7156;
        ChannelMessage t;
        t <- mod_5600.get(16);
        mod_656.put(1, t);
    endrule
    rule rule_7157;
        ChannelMessage t;
        t <- mod_5600.get(39);
        mod_1599.put(1, t);
    endrule
    rule rule_7158;
        ChannelMessage t;
        t <- mod_492.get(0);
        mod_5313.put(115, t);
    endrule
    rule rule_7159;
        ChannelMessage t;
        t <- mod_5166.get(3);
        mod_5646.put(0, t);
    endrule
    rule rule_7160;
        ChannelMessage t;
        t <- mod_5316.get(0);
        mod_533.put(4, t);
    endrule
    rule rule_7161;
        ChannelMessage t;
        t <- mod_5484.get(0);
        mod_779.put(4, t);
    endrule
    rule rule_7162;
        ChannelMessage t;
        t <- mod_5309.get(80);
        mod_3280.put(0, t);
    endrule
    rule rule_7163;
        ChannelMessage t;
        t <- mod_5456.get(0);
        mod_1640.put(2, t);
    endrule
    rule rule_7164;
        ChannelMessage t;
        t <- mod_5442.get(0);
        mod_4592.put(2, t);
    endrule
    rule rule_7165;
        ChannelMessage t;
        t <- mod_3813.get(0);
        mod_5319.put(0, t);
    endrule
    rule rule_7166;
        ChannelMessage t;
        t <- mod_2255.get(0);
        mod_5379.put(0, t);
    endrule
    rule rule_7167;
        ChannelMessage t;
        t <- mod_5309.get(86);
        mod_3526.put(0, t);
    endrule
    rule rule_7168;
        ChannelMessage t;
        t <- mod_2501.get(1);
        mod_5313.put(66, t);
    endrule
    rule rule_7169;
        ChannelMessage t;
        t <- mod_5309.get(30);
        mod_1230.put(0, t);
    endrule
    rule rule_7170;
        ChannelMessage t;
        t <- mod_5439.get(0);
        mod_4346.put(4, t);
    endrule
    rule rule_7171;
        ChannelMessage t;
        t <- mod_5285.get(0);
        mod_861.put(4, t);
    endrule
    rule rule_7172;
        ChannelMessage t;
        t <- mod_410.get(0);
        mod_5267.put(0, t);
    endrule
    rule rule_7173;
        ChannelMessage t;
        t <- mod_5600.get(77);
        mod_3157.put(1, t);
    endrule
    rule rule_7174;
        ChannelMessage t;
        t <- mod_1025.get(0);
        mod_5624.put(0, t);
    endrule
    rule rule_7175;
        ChannelMessage t;
        t <- mod_5607.get(0);
        mod_3690.put(2, t);
    endrule
    rule rule_7176;
        ChannelMessage t;
        t <- mod_5309.get(57);
        mod_2337.put(0, t);
    endrule
    rule rule_7177;
        ChannelMessage t;
        t <- mod_5606.get(0);
        mod_3567.put(3, t);
    endrule
    rule rule_7178;
        ChannelMessage t;
        t <- mod_5520.get(0);
        mod_4346.put(3, t);
    endrule
    rule rule_7179;
        ChannelMessage t;
        t <- mod_3321.get(3);
        mod_5576.put(0, t);
    endrule
    rule rule_7180;
        ChannelMessage t;
        t <- mod_5638.get(0);
        mod_4797.put(2, t);
    endrule
    rule rule_7181;
        ChannelMessage t;
        t <- mod_2296.get(0);
        mod_5313.put(71, t);
    endrule
    rule rule_7182;
        ChannelMessage t;
        t <- mod_2255.get(2);
        mod_5313.put(72, t);
    endrule
    rule rule_7183;
        ChannelMessage t;
        t <- mod_5309.get(88);
        mod_3608.put(0, t);
    endrule
    rule rule_7184;
        ChannelMessage t;
        t <- mod_4059.get(1);
        mod_5313.put(28, t);
    endrule
    rule rule_7185;
        ChannelMessage t;
        t <- mod_2870.get(0);
        mod_5313.put(57, t);
    endrule
    rule rule_7186;
        ChannelMessage t;
        t <- mod_5431.get(0);
        mod_41.put(3, t);
    endrule
    rule rule_7187;
        ChannelMessage t;
        t <- mod_3403.get(2);
        mod_5504.put(0, t);
    endrule
    rule rule_7188;
        ChannelMessage t;
        t <- mod_2993.get(2);
        mod_5258.put(0, t);
    endrule
    rule rule_7189;
        ChannelMessage t;
        t <- mod_205.get(0);
        mod_5341.put(0, t);
    endrule
    rule rule_7190;
        ChannelMessage t;
        t <- mod_5309.get(47);
        mod_1927.put(0, t);
    endrule
    rule rule_7191;
        ChannelMessage t;
        t <- mod_5295.get(0);
        mod_3280.put(2, t);
    endrule
    rule rule_7192;
        ChannelMessage t;
        t <- mod_656.get(3);
        mod_5601.put(0, t);
    endrule
    rule rule_7193;
        ChannelMessage t;
        t <- mod_1066.get(1);
        mod_5554.put(0, t);
    endrule
    rule rule_7194;
        ChannelMessage t;
        t <- mod_533.get(0);
        mod_5557.put(0, t);
    endrule
    rule rule_7195;
        ChannelMessage t;
        t <- mod_5572.get(0);
        mod_943.put(3, t);
    endrule
    rule rule_7196;
        ChannelMessage t;
        t <- mod_5125.get(3);
        mod_5446.put(0, t);
    endrule
    rule rule_7197;
        ChannelMessage t;
        t <- mod_2624.get(0);
        mod_5324.put(0, t);
    endrule
    rule rule_7198;
        ChannelMessage t;
        t <- mod_5309.get(110);
        mod_4510.put(0, t);
    endrule
    rule rule_7199;
        ChannelMessage t;
        t <- mod_5377.get(0);
        mod_5600.put(1, t);
    endrule
    rule rule_7200;
        ChannelMessage t;
        t <- mod_4141.get(0);
        mod_5467.put(0, t);
    endrule
    rule rule_7201;
        ChannelMessage t;
        t <- mod_205.get(2);
        mod_5577.put(0, t);
    endrule
    rule rule_7202;
        ChannelMessage t;
        t <- mod_5309.get(56);
        mod_2296.put(0, t);
    endrule
    rule rule_7203;
        ChannelMessage t;
        t <- mod_3116.get(0);
        mod_5449.put(0, t);
    endrule
    rule rule_7204;
        ChannelMessage t;
        t <- mod_4961.get(0);
        mod_5564.put(0, t);
    endrule
    rule rule_7205;
        ChannelMessage t;
        t <- mod_5486.get(0);
        mod_5043.put(2, t);
    endrule
    rule rule_7206;
        ChannelMessage t;
        t <- mod_3649.get(1);
        mod_5491.put(0, t);
    endrule
    rule rule_7207;
        ChannelMessage t;
        t <- mod_4633.get(0);
        mod_5492.put(0, t);
    endrule
    rule rule_7208;
        ChannelMessage t;
        t <- mod_5441.get(0);
        mod_1845.put(2, t);
    endrule
    rule rule_7209;
        ChannelMessage t;
        t <- mod_5515.get(0);
        mod_2583.put(2, t);
    endrule
    rule rule_7210;
        ChannelMessage t;
        t <- mod_5615.get(0);
        mod_2624.put(3, t);
    endrule
    rule rule_7211;
        ChannelMessage t;
        t <- mod_5368.get(0);
        mod_4510.put(4, t);
    endrule
    rule rule_7212;
        ChannelMessage t;
        t <- mod_3895.get(2);
        mod_5288.put(0, t);
    endrule
    rule rule_7213;
        ChannelMessage t;
        t <- mod_1763.get(0);
        mod_5619.put(0, t);
    endrule
    rule rule_7214;
        ChannelMessage t;
        t <- mod_5521.get(0);
        mod_3649.put(2, t);
    endrule
    rule rule_7215;
        ChannelMessage t;
        t <- mod_5600.get(49);
        mod_2009.put(1, t);
    endrule
    rule rule_7216;
        ChannelMessage t;
        t <- mod_4838.get(2);
        mod_5397.put(0, t);
    endrule
    rule rule_7217;
        ChannelMessage t;
        t <- mod_5434.get(0);
        mod_1107.put(4, t);
    endrule
    rule rule_7218;
        ChannelMessage t;
        t <- mod_5489.get(0);
        mod_164.put(4, t);
    endrule
    rule rule_7219;
        ChannelMessage t;
        t <- mod_2378.get(2);
        mod_5313.put(69, t);
    endrule
    rule rule_7220;
        ChannelMessage t;
        t <- mod_5309.get(33);
        mod_1353.put(0, t);
    endrule
    rule rule_7221;
        ChannelMessage t;
        t <- mod_5372.get(0);
        mod_5326.put(0, t);
    endrule
    rule rule_7222;
        ChannelMessage t;
        t <- mod_5270.get(0);
        mod_2296.put(3, t);
    endrule
    rule rule_7223;
        ChannelMessage t;
        t <- mod_5600.get(14);
        mod_574.put(1, t);
    endrule
    rule rule_7224;
        ChannelMessage t;
        t <- mod_0.get(3);
        mod_5351.put(0, t);
    endrule
    rule rule_7225;
        ChannelMessage t;
        t <- mod_451.get(0);
        mod_5313.put(116, t);
    endrule
    rule rule_7226;
        ChannelMessage t;
        t <- mod_3362.get(0);
        mod_5323.put(0, t);
    endrule
    rule rule_7227;
        ChannelMessage t;
        t <- mod_5309.get(18);
        mod_738.put(0, t);
    endrule
    rule rule_7228;
        ChannelMessage t;
        t <- mod_5328.get(0);
        mod_123.put(2, t);
    endrule
    rule rule_7229;
        ChannelMessage t;
        t <- mod_3198.get(0);
        mod_5448.put(0, t);
    endrule
    rule rule_7230;
        ChannelMessage t;
        t <- mod_4305.get(3);
        mod_5438.put(0, t);
    endrule
    rule rule_7231;
        ChannelMessage t;
        t <- mod_2952.get(3);
        mod_5408.put(0, t);
    endrule
    rule rule_7232;
        ChannelMessage t;
        t <- mod_5309.get(5);
        mod_205.put(0, t);
    endrule
    rule rule_7233;
        ChannelMessage t;
        t <- mod_5309.get(45);
        mod_1845.put(0, t);
    endrule
    rule rule_7234;
        ChannelMessage t;
        t <- mod_5309.get(49);
        mod_2009.put(0, t);
    endrule
    rule rule_7235;
        ChannelMessage t;
        t <- mod_5595.get(0);
        mod_2665.put(4, t);
    endrule
    rule rule_7236;
        ChannelMessage t;
        t <- mod_5600.get(105);
        mod_4305.put(1, t);
    endrule
    rule rule_7237;
        ChannelMessage t;
        t <- mod_369.get(2);
        mod_5452.put(0, t);
    endrule
    rule rule_7238;
        ChannelMessage t;
        t <- mod_615.get(2);
        mod_5313.put(112, t);
    endrule
    rule rule_7239;
        ChannelMessage t;
        t <- mod_2009.get(1);
        mod_5321.put(0, t);
    endrule
    rule rule_7240;
        ChannelMessage t;
        t <- mod_5359.get(0);
        mod_205.put(3, t);
    endrule
    rule rule_7241;
        ChannelMessage t;
        t <- mod_5600.get(126);
        mod_5166.put(1, t);
    endrule
    rule rule_7242;
        ChannelMessage t;
        t <- mod_5309.get(16);
        mod_656.put(0, t);
    endrule
    rule rule_7243;
        ChannelMessage t;
        t <- mod_1271.get(3);
        mod_5313.put(96, t);
    endrule
    rule rule_7244;
        ChannelMessage t;
        t <- mod_2050.get(1);
        mod_5325.put(0, t);
    endrule
    rule rule_7245;
        ChannelMessage t;
        t <- mod_5504.get(0);
        mod_3403.put(3, t);
    endrule
    rule rule_7246;
        ChannelMessage t;
        t <- mod_123.get(2);
        mod_5358.put(0, t);
    endrule
    rule rule_7247;
        ChannelMessage t;
        t <- mod_5575.get(0);
        mod_2624.put(4, t);
    endrule
    rule rule_7248;
        ChannelMessage t;
        t <- mod_5271.get(0);
        mod_1681.put(4, t);
    endrule
    rule rule_7249;
        ChannelMessage t;
        t <- mod_2337.get(0);
        mod_5421.put(0, t);
    endrule
    rule rule_7250;
        ChannelMessage t;
        t <- mod_4551.get(3);
        mod_5313.put(16, t);
    endrule
    rule rule_7251;
        ChannelMessage t;
        t <- mod_5309.get(34);
        mod_1394.put(0, t);
    endrule
    rule rule_7252;
        ChannelMessage t;
        t <- mod_5363.get(0);
        mod_2501.put(4, t);
    endrule
    rule rule_7253;
        ChannelMessage t;
        t <- mod_5480.get(0);
        mod_451.put(3, t);
    endrule
    rule rule_7254;
        ChannelMessage t;
        t <- mod_1066.get(3);
        mod_5262.put(0, t);
    endrule
    rule rule_7255;
        ChannelMessage t;
        t <- mod_5309.get(89);
        mod_3649.put(0, t);
    endrule
    rule rule_7256;
        ChannelMessage t;
        t <- mod_5542.get(0);
        mod_1886.put(3, t);
    endrule
    rule rule_7257;
        ChannelMessage t;
        t <- mod_287.get(2);
        mod_5394.put(0, t);
    endrule
    rule rule_7258;
        ChannelMessage t;
        t <- mod_1968.get(3);
        mod_5261.put(0, t);
    endrule
    rule rule_7259;
        ChannelMessage t;
        t <- mod_5647.get(0);
        mod_3157.put(2, t);
    endrule
    rule rule_7260;
        ChannelMessage t;
        t <- mod_5600.get(9);
        mod_369.put(1, t);
    endrule
    rule rule_7261;
        ChannelMessage t;
        t <- mod_5613.get(0);
        mod_4879.put(3, t);
    endrule
    rule rule_7262;
        ChannelMessage t;
        t <- mod_2173.get(0);
        mod_5573.put(0, t);
    endrule
    rule rule_7263;
        ChannelMessage t;
        t <- mod_2173.get(1);
        mod_5510.put(0, t);
    endrule
    rule rule_7264;
        ChannelMessage t;
        t <- mod_5639.get(0);
        mod_779.put(3, t);
    endrule
    rule rule_7265;
        ChannelMessage t;
        t <- mod_5309.get(96);
        mod_3936.put(0, t);
    endrule
    rule rule_7266;
        ChannelMessage t;
        t <- mod_5556.get(0);
        mod_3280.put(3, t);
    endrule
    rule rule_7267;
        ChannelMessage t;
        t <- mod_4305.get(0);
        mod_5594.put(0, t);
    endrule
    rule rule_7268;
        ChannelMessage t;
        t <- mod_246.get(0);
        mod_5337.put(0, t);
    endrule
    rule rule_7269;
        ChannelMessage t;
        t <- mod_4469.get(3);
        mod_5275.put(0, t);
    endrule
    rule rule_7270;
        ChannelMessage t;
        t <- mod_5506.get(0);
        mod_3854.put(3, t);
    endrule
    rule rule_7271;
        ChannelMessage t;
        t <- mod_5427.get(0);
        mod_4592.put(3, t);
    endrule
    rule rule_7272;
        ChannelMessage t;
        t <- mod_5600.get(122);
        mod_5002.put(1, t);
    endrule
    rule rule_7273;
        ChannelMessage t;
        t <- mod_5309.get(26);
        mod_1066.put(0, t);
    endrule
    rule rule_7274;
        ChannelMessage t;
        t <- mod_1927.get(3);
        mod_5349.put(0, t);
    endrule
    rule rule_7275;
        ChannelMessage t;
        t <- mod_5617.get(0);
        mod_1476.put(3, t);
    endrule
    rule rule_7276;
        ChannelMessage t;
        t <- mod_2788.get(3);
        mod_5273.put(0, t);
    endrule
    rule rule_7277;
        ChannelMessage t;
        t <- mod_5309.get(119);
        mod_4879.put(0, t);
    endrule
    rule rule_7278;
        ChannelMessage t;
        t <- mod_4674.get(2);
        mod_5320.put(0, t);
    endrule
    rule rule_7279;
        ChannelMessage t;
        t <- mod_5309.get(9);
        mod_369.put(0, t);
    endrule
    rule rule_7280;
        ChannelMessage t;
        t <- mod_4264.get(1);
        mod_5437.put(0, t);
    endrule
    rule rule_7281;
        ChannelMessage t;
        t <- mod_3608.get(1);
        mod_5313.put(39, t);
    endrule
    rule rule_7282;
        ChannelMessage t;
        t <- mod_5269.get(0);
        mod_1558.put(3, t);
    endrule
    rule rule_7283;
        ChannelMessage t;
        t <- mod_5537.get(0);
        mod_2419.put(3, t);
    endrule
    rule rule_7284;
        ChannelMessage t;
        t <- mod_1394.get(0);
        mod_5313.put(93, t);
    endrule
    rule rule_7285;
        ChannelMessage t;
        t <- mod_5633.get(0);
        mod_4428.put(2, t);
    endrule
    rule rule_7286;
        ChannelMessage t;
        t <- mod_82.get(2);
        mod_5445.put(0, t);
    endrule
    rule rule_7287;
        ChannelMessage t;
        t <- mod_1353.get(3);
        mod_5313.put(94, t);
    endrule
    rule rule_7288;
        ChannelMessage t;
        t <- mod_5309.get(116);
        mod_4756.put(0, t);
    endrule
    rule rule_7289;
        ChannelMessage t;
        t <- mod_3690.get(1);
        mod_5402.put(0, t);
    endrule
    rule rule_7290;
        ChannelMessage t;
        t <- mod_5600.get(127);
        mod_5207.put(1, t);
    endrule
    rule rule_7291;
        ChannelMessage t;
        t <- mod_5388.get(0);
        mod_5002.put(2, t);
    endrule
    rule rule_7292;
        ChannelMessage t;
        t <- mod_4715.get(2);
        mod_5317.put(0, t);
    endrule
    rule rule_7293;
        ChannelMessage t;
        t <- mod_5432.get(0);
        mod_5166.put(2, t);
    endrule
    rule rule_7294;
        ChannelMessage t;
        t <- mod_1968.get(2);
        mod_5538.put(0, t);
    endrule
    rule rule_7295;
        ChannelMessage t;
        t <- mod_3772.get(2);
        mod_5430.put(0, t);
    endrule
    rule rule_7296;
        ChannelMessage t;
        t <- mod_5418.get(0);
        mod_5084.put(4, t);
    endrule
    rule rule_7297;
        ChannelMessage t;
        t <- mod_5600.get(119);
        mod_4879.put(1, t);
    endrule
    rule rule_7298;
        ChannelMessage t;
        t <- mod_1148.get(3);
        mod_5597.put(0, t);
    endrule
    rule rule_7299;
        ChannelMessage t;
        t <- mod_2829.get(1);
        mod_5313.put(58, t);
    endrule
    rule rule_7300;
        ChannelMessage t;
        t <- mod_5351.get(0);
        mod_0.put(3, t);
    endrule
    rule rule_7301;
        ChannelMessage t;
        t <- mod_5360.get(0);
        mod_246.put(4, t);
    endrule
    rule rule_7302;
        ChannelMessage t;
        t <- mod_5600.get(85);
        mod_3485.put(1, t);
    endrule
    rule rule_7303;
        ChannelMessage t;
        t <- mod_5409.get(0);
        mod_1763.put(4, t);
    endrule
    rule rule_7304;
        ChannelMessage t;
        t <- mod_5309.get(44);
        mod_1804.put(0, t);
    endrule
    rule rule_7305;
        ChannelMessage t;
        t <- mod_5449.get(0);
        mod_3116.put(3, t);
    endrule
    rule rule_7306;
        ChannelMessage t;
        t <- mod_4264.get(3);
        mod_5336.put(0, t);
    endrule
    rule rule_7307;
        ChannelMessage t;
        t <- mod_4387.get(1);
        mod_5313.put(20, t);
    endrule
    rule rule_7308;
        ChannelMessage t;
        t <- mod_3895.get(0);
        mod_5259.put(0, t);
    endrule
    rule rule_7309;
        ChannelMessage t;
        t <- mod_5600.get(2);
        mod_82.put(1, t);
    endrule
    rule rule_7310;
        ChannelMessage t;
        t <- mod_5309.get(68);
        mod_2788.put(0, t);
    endrule
    rule rule_7311;
        ChannelMessage t;
        t <- mod_1107.get(3);
        mod_5332.put(0, t);
    endrule
    rule rule_7312;
        ChannelMessage t;
        t <- mod_1640.get(3);
        mod_5282.put(0, t);
    endrule
    rule rule_7313;
        ChannelMessage t;
        t <- mod_5305.get(0);
        mod_1927.put(2, t);
    endrule
    rule rule_7314;
        ChannelMessage t;
        t <- mod_5438.get(0);
        mod_4305.put(3, t);
    endrule
    rule rule_7315;
        ChannelMessage t;
        t <- mod_5474.get(0);
        mod_615.put(3, t);
    endrule
    rule rule_7316;
        ChannelMessage t;
        t <- mod_41.get(0);
        mod_5407.put(0, t);
    endrule
    rule rule_7317;
        ChannelMessage t;
        t <- mod_2788.get(2);
        mod_5503.put(0, t);
    endrule
    rule rule_7318;
        ChannelMessage t;
        t <- mod_5395.get(0);
        mod_5207.put(2, t);
    endrule
    rule rule_7319;
        ChannelMessage t;
        t <- mod_5389.get(0);
        mod_4264.put(2, t);
    endrule
    rule rule_7320;
        ChannelMessage t;
        t <- mod_5256.get(0);
        mod_3936.put(4, t);
    endrule
    rule rule_7321;
        ChannelMessage t;
        t <- mod_5497.get(0);
        mod_2460.put(3, t);
    endrule
    rule rule_7322;
        ChannelMessage t;
        t <- mod_697.get(0);
        mod_5561.put(0, t);
    endrule
    rule rule_7323;
        ChannelMessage t;
        t <- mod_1148.get(2);
        mod_5644.put(0, t);
    endrule
    rule rule_7324;
        ChannelMessage t;
        t <- mod_5600.get(24);
        mod_984.put(1, t);
    endrule
    rule rule_7325;
        ChannelMessage t;
        t <- mod_4223.get(2);
        mod_5313.put(24, t);
    endrule
    rule rule_7326;
        ChannelMessage t;
        t <- mod_1804.get(2);
        mod_5348.put(0, t);
    endrule
    rule rule_7327;
        ChannelMessage t;
        t <- mod_4182.get(2);
        mod_5313.put(25, t);
    endrule
    rule rule_7328;
        ChannelMessage t;
        t <- mod_1640.get(1);
        mod_5456.put(0, t);
    endrule
    rule rule_7329;
        ChannelMessage t;
        t <- mod_5309.get(109);
        mod_4469.put(0, t);
    endrule
    rule rule_7330;
        ChannelMessage t;
        t <- mod_4018.get(0);
        mod_5289.put(0, t);
    endrule
    rule rule_7331;
        ChannelMessage t;
        t <- mod_5600.get(10);
        mod_410.put(1, t);
    endrule
    rule rule_7332;
        ChannelMessage t;
        t <- mod_3157.get(1);
        mod_5266.put(0, t);
    endrule
    rule rule_7333;
        ChannelMessage t;
        t <- mod_5353.get(0);
        mod_984.put(3, t);
    endrule
    rule rule_7334;
        ChannelMessage t;
        t <- mod_3321.get(2);
        mod_5281.put(0, t);
    endrule
    rule rule_7335;
        ChannelMessage t;
        t <- mod_4633.get(2);
        mod_5565.put(0, t);
    endrule
    rule rule_7336;
        ChannelMessage t;
        t <- mod_2583.get(2);
        mod_5293.put(0, t);
    endrule
    rule rule_7337;
        ChannelMessage t;
        t <- mod_1271.get(1);
        mod_5301.put(0, t);
    endrule
    rule rule_7338;
        ChannelMessage t;
        t <- mod_5290.get(0);
        mod_1763.put(3, t);
    endrule
    rule rule_7339;
        ChannelMessage t;
        t <- mod_5482.get(0);
        mod_1394.put(4, t);
    endrule
    rule rule_7340;
        ChannelMessage t;
        t <- mod_4387.get(2);
        mod_5525.put(0, t);
    endrule
    rule rule_7341;
        ChannelMessage t;
        t <- mod_5550.get(0);
        mod_451.put(2, t);
    endrule
    rule rule_7342;
        ChannelMessage t;
        t <- mod_5600.get(63);
        mod_2583.put(1, t);
    endrule
    rule rule_7343;
        ChannelMessage t;
        t <- mod_5526.get(0);
        mod_5309.put(1, t);
    endrule
    rule rule_7344;
        ChannelMessage t;
        t <- mod_5600.get(65);
        mod_2665.put(1, t);
    endrule
    rule rule_7345;
        ChannelMessage t;
        t <- mod_2911.get(2);
        mod_5333.put(0, t);
    endrule
    rule rule_7346;
        ChannelMessage t;
        t <- mod_5309.get(97);
        mod_3977.put(0, t);
    endrule
    rule rule_7347;
        ChannelMessage t;
        t <- mod_5379.get(0);
        mod_2255.put(4, t);
    endrule
    rule rule_7348;
        ChannelMessage t;
        t <- mod_5560.get(0);
        mod_4059.put(3, t);
    endrule
    rule rule_7349;
        ChannelMessage t;
        t <- mod_5600.get(53);
        mod_2173.put(1, t);
    endrule
    rule rule_7350;
        ChannelMessage t;
        t <- mod_1804.get(3);
        mod_5628.put(0, t);
    endrule
    rule rule_7351;
        ChannelMessage t;
        t <- mod_2173.get(3);
        mod_5313.put(74, t);
    endrule
    rule rule_7352;
        ChannelMessage t;
        t <- mod_1845.get(3);
        mod_5313.put(82, t);
    endrule
    rule rule_7353;
        ChannelMessage t;
        t <- mod_5485.get(0);
        mod_2747.put(4, t);
    endrule
    rule rule_7354;
        ChannelMessage t;
        t <- mod_4018.get(2);
        mod_5313.put(29, t);
    endrule
    rule rule_7355;
        ChannelMessage t;
        t <- mod_5333.get(0);
        mod_2911.put(4, t);
    endrule
    rule rule_7356;
        ChannelMessage t;
        t <- mod_5347.get(0);
        mod_656.put(4, t);
    endrule
    rule rule_7357;
        ChannelMessage t;
        t <- mod_4756.get(0);
        mod_5265.put(0, t);
    endrule
    rule rule_7358;
        ChannelMessage t;
        t <- mod_5600.get(89);
        mod_3649.put(1, t);
    endrule
    rule rule_7359;
        ChannelMessage t;
        t <- mod_5561.get(0);
        mod_697.put(3, t);
    endrule
    rule rule_7360;
        ChannelMessage t;
        t <- mod_1107.get(0);
        mod_5313.put(100, t);
    endrule
    rule rule_7361;
        ChannelMessage t;
        t <- mod_5166.get(0);
        mod_5432.put(0, t);
    endrule
    rule rule_7362;
        ChannelMessage t;
        t <- mod_2665.get(2);
        mod_5249.put(0, t);
    endrule
    rule rule_7363;
        ChannelMessage t;
        t <- mod_5544.get(0);
        mod_3895.put(4, t);
    endrule
    rule rule_7364;
        ChannelMessage t;
        t <- mod_5563.get(0);
        mod_2255.put(2, t);
    endrule
    rule rule_7365;
        ChannelMessage t;
        t <- mod_5309.get(77);
        mod_3157.put(0, t);
    endrule
    rule rule_7366;
        ChannelMessage t;
        t <- mod_5309.get(122);
        mod_5002.put(0, t);
    endrule
    rule rule_7367;
        ChannelMessage t;
        t <- mod_5381.get(0);
        mod_738.put(2, t);
    endrule
    rule rule_7368;
        ChannelMessage t;
        t <- mod_1476.get(0);
        mod_5414.put(0, t);
    endrule
    rule rule_7369;
        ChannelMessage t;
        t <- mod_5600.get(45);
        mod_1845.put(1, t);
    endrule
    rule rule_7370;
        ChannelMessage t;
        t <- mod_533.get(2);
        mod_5488.put(0, t);
    endrule
    rule rule_7371;
        ChannelMessage t;
        t <- mod_4141.get(3);
        mod_5313.put(26, t);
    endrule
    rule rule_7372;
        ChannelMessage t;
        t <- mod_3526.get(0);
        mod_5313.put(41, t);
    endrule
    rule rule_7373;
        ChannelMessage t;
        t <- mod_5293.get(0);
        mod_2583.put(3, t);
    endrule
    rule rule_7374;
        ChannelMessage t;
        t <- mod_2952.get(1);
        mod_5313.put(55, t);
    endrule
    rule rule_7375;
        ChannelMessage t;
        t <- mod_5423.get(0);
        mod_1025.put(4, t);
    endrule
    rule rule_7376;
        ChannelMessage t;
        t <- mod_5411.get(0);
        mod_1845.put(3, t);
    endrule
    rule rule_7377;
        ChannelMessage t;
        t <- mod_5382.get(0);
        mod_902.put(3, t);
    endrule
    rule rule_7378;
        ChannelMessage t;
        t <- mod_5286.get(0);
        mod_2542.put(3, t);
    endrule
    rule rule_7379;
        ChannelMessage t;
        t <- mod_5600.get(43);
        mod_1763.put(1, t);
    endrule
    rule rule_7380;
        ChannelMessage t;
        t <- mod_2296.get(2);
        mod_5551.put(0, t);
    endrule
    rule rule_7381;
        ChannelMessage t;
        t <- mod_5436.get(0);
        mod_820.put(2, t);
    endrule
    rule rule_7382;
        ChannelMessage t;
        t <- mod_1394.get(1);
        mod_5482.put(0, t);
    endrule
    rule rule_7383;
        ChannelMessage t;
        t <- mod_5361.get(0);
        mod_3813.put(3, t);
    endrule
    rule rule_7384;
        ChannelMessage t;
        t <- mod_2993.get(0);
        mod_5415.put(0, t);
    endrule
    rule rule_7385;
        ChannelMessage t;
        t <- mod_2460.get(0);
        mod_5497.put(0, t);
    endrule
    rule rule_7386;
        ChannelMessage t;
        t <- mod_246.get(2);
        mod_5360.put(0, t);
    endrule
    rule rule_7387;
        ChannelMessage t;
        t <- mod_1230.get(0);
        mod_5390.put(0, t);
    endrule
    rule rule_7388;
        ChannelMessage t;
        t <- mod_2091.get(1);
        mod_5453.put(0, t);
    endrule
    rule rule_7389;
        ChannelMessage t;
        t <- mod_4838.get(1);
        mod_5458.put(0, t);
    endrule
    rule rule_7390;
        ChannelMessage t;
        t <- mod_5313.get(0);
        mod_5372.put(0, t);
    endrule
    rule rule_7391;
        ChannelMessage t;
        t <- mod_5600.get(19);
        mod_779.put(1, t);
    endrule
    rule rule_7392;
        ChannelMessage t;
        t <- mod_5325.get(0);
        mod_2050.put(4, t);
    endrule
    rule rule_7393;
        ChannelMessage t;
        t <- mod_3444.get(2);
        mod_5508.put(0, t);
    endrule
    rule rule_7394;
        ChannelMessage t;
        t <- mod_2993.get(1);
        mod_5313.put(54, t);
    endrule
    rule rule_7395;
        ChannelMessage t;
        t <- mod_5326.get(0);
        mod_5326.put(1, t);
    endrule
    rule rule_7396;
        ChannelMessage t;
        t <- mod_5437.get(0);
        mod_4264.put(3, t);
    endrule
    rule rule_7397;
        ChannelMessage t;
        t <- mod_5530.get(0);
        mod_1230.put(2, t);
    endrule
    rule rule_7398;
        ChannelMessage t;
        t <- mod_5592.get(0);
        mod_1394.put(2, t);
    endrule
    rule rule_7399;
        ChannelMessage t;
        t <- mod_5600.get(79);
        mod_3239.put(1, t);
    endrule
    rule rule_7400;
        ChannelMessage t;
        t <- mod_5602.get(0);
        mod_1886.put(2, t);
    endrule
    rule rule_7401;
        ChannelMessage t;
        t <- mod_902.get(2);
        mod_5419.put(0, t);
    endrule
    rule rule_7402;
        ChannelMessage t;
        t <- mod_5631.get(0);
        mod_0.put(2, t);
    endrule
    rule rule_7403;
        ChannelMessage t;
        t <- mod_5249.get(0);
        mod_2665.put(2, t);
    endrule
    rule rule_7404;
        ChannelMessage t;
        t <- mod_5600.get(5);
        mod_205.put(1, t);
    endrule
    rule rule_7405;
        ChannelMessage t;
        t <- mod_738.get(3);
        mod_5313.put(109, t);
    endrule
    rule rule_7406;
        ChannelMessage t;
        t <- mod_5309.get(38);
        mod_1558.put(0, t);
    endrule
    rule rule_7407;
        ChannelMessage t;
        t <- mod_5421.get(0);
        mod_2337.put(4, t);
    endrule
    rule rule_7408;
        ChannelMessage t;
        t <- mod_2542.get(2);
        mod_5540.put(0, t);
    endrule
    rule rule_7409;
        ChannelMessage t;
        t <- mod_5348.get(0);
        mod_1804.put(2, t);
    endrule
    rule rule_7410;
        ChannelMessage t;
        t <- mod_5433.get(0);
        mod_861.put(3, t);
    endrule
    rule rule_7411;
        ChannelMessage t;
        t <- mod_4182.get(0);
        mod_5327.put(0, t);
    endrule
    rule rule_7412;
        ChannelMessage t;
        t <- mod_1271.get(2);
        mod_5331.put(0, t);
    endrule
    rule rule_7413;
        ChannelMessage t;
        t <- mod_5330.get(0);
        mod_2378.put(2, t);
    endrule
    rule rule_7414;
        ChannelMessage t;
        t <- mod_615.get(1);
        mod_5479.put(0, t);
    endrule
    rule rule_7415;
        ChannelMessage t;
        t <- mod_2091.get(3);
        mod_5403.put(0, t);
    endrule
    rule rule_7416;
        ChannelMessage t;
        t <- mod_5625.get(0);
        mod_3977.put(4, t);
    endrule
    rule rule_7417;
        ChannelMessage t;
        t <- mod_5350.get(0);
        mod_5377.put(0, t);
    endrule
    rule rule_7418;
        ChannelMessage t;
        t <- mod_820.get(0);
        mod_5436.put(0, t);
    endrule
    rule rule_7419;
        ChannelMessage t;
        t <- mod_738.get(2);
        mod_5362.put(0, t);
    endrule
    rule rule_7420;
        ChannelMessage t;
        t <- mod_1025.get(2);
        mod_5451.put(0, t);
    endrule
    rule rule_7421;
        ChannelMessage t;
        t <- mod_2378.get(0);
        mod_5365.put(0, t);
    endrule
    rule rule_7422;
        ChannelMessage t;
        t <- mod_2829.get(0);
        mod_5608.put(0, t);
    endrule
    rule rule_7423;
        ChannelMessage t;
        t <- mod_5309.get(6);
        mod_246.put(0, t);
    endrule
    rule rule_7424;
        ChannelMessage t;
        t <- mod_5251.get(0);
        mod_328.put(4, t);
    endrule
    rule rule_7425;
        ChannelMessage t;
        t <- mod_4551.get(1);
        mod_5559.put(0, t);
    endrule
    rule rule_7426;
        ChannelMessage t;
        t <- mod_779.get(1);
        mod_5428.put(0, t);
    endrule
    rule rule_7427;
        ChannelMessage t;
        t <- mod_5309.get(58);
        mod_2378.put(0, t);
    endrule
    rule rule_7428;
        ChannelMessage t;
        t <- mod_5600.get(52);
        mod_2132.put(1, t);
    endrule
    rule rule_7429;
        ChannelMessage t;
        t <- mod_5611.get(0);
        mod_1722.put(4, t);
    endrule
    rule rule_7430;
        ChannelMessage t;
        t <- mod_3567.get(1);
        mod_5313.put(40, t);
    endrule
    rule rule_7431;
        ChannelMessage t;
        t <- mod_0.get(1);
        mod_5631.put(0, t);
    endrule
    rule rule_7432;
        ChannelMessage t;
        t <- mod_2583.get(3);
        mod_5515.put(0, t);
    endrule
    rule rule_7433;
        ChannelMessage t;
        t <- mod_5268.get(0);
        mod_2706.put(3, t);
    endrule
    rule rule_7434;
        ChannelMessage t;
        t <- mod_5265.get(0);
        mod_4756.put(3, t);
    endrule
    rule rule_7435;
        ChannelMessage t;
        t <- mod_2419.get(3);
        mod_5313.put(68, t);
    endrule
    rule rule_7436;
        ChannelMessage t;
        t <- mod_2583.get(1);
        mod_5516.put(0, t);
    endrule
    rule rule_7437;
        ChannelMessage t;
        t <- mod_5258.get(0);
        mod_2993.put(4, t);
    endrule
    rule rule_7438;
        ChannelMessage t;
        t <- mod_3403.get(3);
        mod_5596.put(0, t);
    endrule
    rule rule_7439;
        ChannelMessage t;
        t <- mod_5300.get(0);
        mod_4469.put(3, t);
    endrule
    rule rule_7440;
        ChannelMessage t;
        t <- mod_2050.get(2);
        mod_5313.put(77, t);
    endrule
    rule rule_7441;
        ChannelMessage t;
        t <- mod_5539.get(0);
        mod_4592.put(4, t);
    endrule
    rule rule_7442;
        ChannelMessage t;
        t <- mod_2665.get(3);
        mod_5374.put(0, t);
    endrule
    rule rule_7443;
        ChannelMessage t;
        t <- mod_3485.get(2);
        mod_5313.put(42, t);
    endrule
    rule rule_7444;
        ChannelMessage t;
        t <- mod_5466.get(0);
        mod_3075.put(4, t);
    endrule
    rule rule_7445;
        ChannelMessage t;
        t <- mod_5519.get(0);
        mod_4018.put(3, t);
    endrule
    rule rule_7446;
        ChannelMessage t;
        t <- mod_5535.get(0);
        mod_1517.put(2, t);
    endrule
    rule rule_7447;
        ChannelMessage t;
        t <- mod_5407.get(0);
        mod_41.put(2, t);
    endrule
    rule rule_7448;
        ChannelMessage t;
        t <- mod_5450.get(0);
        mod_1722.put(3, t);
    endrule
    rule rule_7449;
        ChannelMessage t;
        t <- mod_5386.get(0);
        mod_1271.put(3, t);
    endrule
    rule rule_7450;
        ChannelMessage t;
        t <- mod_5629.get(0);
        mod_2870.put(2, t);
    endrule
    rule rule_7451;
        ChannelMessage t;
        t <- mod_205.get(1);
        mod_5313.put(122, t);
    endrule
    rule rule_7452;
        ChannelMessage t;
        t <- mod_2337.get(3);
        mod_5502.put(0, t);
    endrule
    rule rule_7453;
        ChannelMessage t;
        t <- mod_4920.get(0);
        mod_5313.put(7, t);
    endrule
    rule rule_7454;
        ChannelMessage t;
        t <- mod_5309.get(71);
        mod_2911.put(0, t);
    endrule
    rule rule_7455;
        ChannelMessage t;
        t <- mod_5493.get(0);
        mod_3977.put(2, t);
    endrule
    rule rule_7456;
        ChannelMessage t;
        t <- mod_82.get(0);
        mod_5313.put(125, t);
    endrule
    rule rule_7457;
        ChannelMessage t;
        t <- mod_5261.get(0);
        mod_1968.put(2, t);
    endrule
    rule rule_7458;
        ChannelMessage t;
        t <- mod_5299.get(0);
        mod_1107.put(2, t);
    endrule
    rule rule_7459;
        ChannelMessage t;
        t <- mod_5309.get(51);
        mod_2091.put(0, t);
    endrule
    rule rule_7460;
        ChannelMessage t;
        t <- mod_5508.get(0);
        mod_3444.put(2, t);
    endrule
    rule rule_7461;
        ChannelMessage t;
        t <- mod_4551.get(2);
        mod_5391.put(0, t);
    endrule
    rule rule_7462;
        ChannelMessage t;
        t <- mod_3977.get(2);
        mod_5478.put(0, t);
    endrule
    rule rule_7463;
        ChannelMessage t;
        t <- mod_5574.get(0);
        mod_4059.put(4, t);
    endrule
    rule rule_7464;
        ChannelMessage t;
        t <- mod_5084.get(3);
        mod_5529.put(0, t);
    endrule
    rule rule_7465;
        ChannelMessage t;
        t <- mod_2542.get(3);
        mod_5313.put(65, t);
    endrule
    rule rule_7466;
        ChannelMessage t;
        t <- mod_4018.get(3);
        mod_5519.put(0, t);
    endrule
    rule rule_7467;
        ChannelMessage t;
        t <- mod_328.get(0);
        mod_5548.put(0, t);
    endrule
    rule rule_7468;
        ChannelMessage t;
        t <- mod_4059.get(0);
        mod_5574.put(0, t);
    endrule
    rule rule_7469;
        ChannelMessage t;
        t <- mod_5309.get(92);
        mod_3772.put(0, t);
    endrule
    rule rule_7470;
        ChannelMessage t;
        t <- mod_5324.get(0);
        mod_2624.put(2, t);
    endrule
    rule rule_7471;
        ChannelMessage t;
        t <- mod_5499.get(0);
        mod_4100.put(3, t);
    endrule
    rule rule_7472;
        ChannelMessage t;
        t <- mod_1845.get(0);
        mod_5329.put(0, t);
    endrule
    rule rule_7473;
        ChannelMessage t;
        t <- mod_2132.get(0);
        mod_5571.put(0, t);
    endrule
    rule rule_7474;
        ChannelMessage t;
        t <- mod_5207.get(1);
        mod_5395.put(0, t);
    endrule
    rule rule_7475;
        ChannelMessage t;
        t <- mod_5309.get(17);
        mod_697.put(0, t);
    endrule
    rule rule_7476;
        ChannelMessage t;
        t <- mod_5339.get(0);
        mod_820.put(4, t);
    endrule
    rule rule_7477;
        ChannelMessage t;
        t <- mod_2952.get(2);
        mod_5514.put(0, t);
    endrule
    rule rule_7478;
        ChannelMessage t;
        t <- mod_5349.get(0);
        mod_1927.put(3, t);
    endrule
    rule rule_7479;
        ChannelMessage t;
        t <- mod_5533.get(0);
        mod_2132.put(3, t);
    endrule
    rule rule_7480;
        ChannelMessage t;
        t <- mod_4141.get(2);
        mod_5425.put(0, t);
    endrule
    rule rule_7481;
        ChannelMessage t;
        t <- mod_4879.get(1);
        mod_5622.put(0, t);
    endrule
    rule rule_7482;
        ChannelMessage t;
        t <- mod_5582.get(0);
        mod_1968.put(4, t);
    endrule
    rule rule_7483;
        ChannelMessage t;
        t <- mod_4305.get(1);
        mod_5413.put(0, t);
    endrule
    rule rule_7484;
        ChannelMessage t;
        t <- mod_5084.get(0);
        mod_5614.put(0, t);
    endrule
    rule rule_7485;
        ChannelMessage t;
        t <- mod_5568.get(0);
        mod_1681.put(2, t);
    endrule
    rule rule_7486;
        ChannelMessage t;
        t <- mod_5503.get(0);
        mod_2788.put(3, t);
    endrule
    rule rule_7487;
        ChannelMessage t;
        t <- mod_1681.get(1);
        mod_5271.put(0, t);
    endrule
    rule rule_7488;
        ChannelMessage t;
        t <- mod_5253.get(0);
        mod_5043.put(3, t);
    endrule
    rule rule_7489;
        ChannelMessage t;
        t <- mod_4223.get(1);
        mod_5511.put(0, t);
    endrule
    rule rule_7490;
        ChannelMessage t;
        t <- mod_5373.get(0);
        mod_4715.put(2, t);
    endrule
    rule rule_7491;
        ChannelMessage t;
        t <- mod_5404.get(0);
        mod_492.put(2, t);
    endrule
    rule rule_7492;
        ChannelMessage t;
        t <- mod_3936.get(2);
        mod_5313.put(31, t);
    endrule
    rule rule_7493;
        ChannelMessage t;
        t <- mod_5600.get(25);
        mod_1025.put(1, t);
    endrule
    rule rule_7494;
        ChannelMessage t;
        t <- mod_1312.get(1);
        mod_5304.put(0, t);
    endrule
    rule rule_7495;
        ChannelMessage t;
        t <- mod_164.get(1);
        mod_5313.put(123, t);
    endrule
    rule rule_7496;
        ChannelMessage t;
        t <- mod_2583.get(0);
        mod_5313.put(64, t);
    endrule
    rule rule_7497;
        ChannelMessage t;
        t <- mod_3034.get(2);
        mod_5637.put(0, t);
    endrule
    rule rule_7498;
        ChannelMessage t;
        t <- mod_5309.get(83);
        mod_3403.put(0, t);
    endrule
    rule rule_7499;
        ChannelMessage t;
        t <- mod_5435.get(0);
        mod_2870.put(4, t);
    endrule
    rule rule_7500;
        ChannelMessage t;
        t <- mod_3690.get(2);
        mod_5313.put(37, t);
    endrule
    rule rule_7501;
        ChannelMessage t;
        t <- mod_5376.get(0);
        mod_4469.put(2, t);
    endrule
    rule rule_7502;
        ChannelMessage t;
        t <- mod_5309.get(40);
        mod_1640.put(0, t);
    endrule
    rule rule_7503;
        ChannelMessage t;
        t <- mod_5494.get(0);
        mod_3444.put(3, t);
    endrule
    rule rule_7504;
        ChannelMessage t;
        t <- mod_5567.get(0);
        mod_4715.put(4, t);
    endrule
    rule rule_7505;
        ChannelMessage t;
        t <- mod_5600.get(61);
        mod_2501.put(1, t);
    endrule
    rule rule_7506;
        ChannelMessage t;
        t <- mod_4674.get(1);
        mod_5313.put(13, t);
    endrule
    rule rule_7507;
        ChannelMessage t;
        t <- mod_2460.get(3);
        mod_5648.put(0, t);
    endrule
    rule rule_7508;
        ChannelMessage t;
        t <- mod_1517.get(2);
        mod_5584.put(0, t);
    endrule
    rule rule_7509;
        ChannelMessage t;
        t <- mod_5600.get(12);
        mod_492.put(1, t);
    endrule
    rule rule_7510;
        ChannelMessage t;
        t <- mod_2706.get(0);
        mod_5313.put(61, t);
    endrule
    rule rule_7511;
        ChannelMessage t;
        t <- mod_5569.get(0);
        mod_2091.put(3, t);
    endrule
    rule rule_7512;
        ChannelMessage t;
        t <- mod_5309.get(42);
        mod_1722.put(0, t);
    endrule
    rule rule_7513;
        ChannelMessage t;
        t <- mod_5416.get(0);
        mod_2214.put(3, t);
    endrule
    rule rule_7514;
        ChannelMessage t;
        t <- mod_5614.get(0);
        mod_5084.put(2, t);
    endrule
    rule rule_7515;
        ChannelMessage t;
        t <- mod_5642.get(0);
        mod_3731.put(2, t);
    endrule
    rule rule_7516;
        ChannelMessage t;
        t <- mod_5344.get(0);
        mod_5248.put(0, t);
    endrule
    rule rule_7517;
        ChannelMessage t;
        t <- mod_5507.get(0);
        mod_3198.put(3, t);
    endrule
    rule rule_7518;
        ChannelMessage t;
        t <- mod_492.get(3);
        mod_5610.put(0, t);
    endrule
    rule rule_7519;
        ChannelMessage t;
        t <- mod_5002.get(3);
        mod_5552.put(0, t);
    endrule
    rule rule_7520;
        ChannelMessage t;
        t <- mod_5250.get(0);
        mod_4428.put(4, t);
    endrule
    rule rule_7521;
        ChannelMessage t;
        t <- mod_943.get(0);
        mod_5334.put(0, t);
    endrule
    rule rule_7522;
        ChannelMessage t;
        t <- mod_1558.get(1);
        mod_5313.put(89, t);
    endrule
    rule rule_7523;
        ChannelMessage t;
        t <- mod_1845.get(1);
        mod_5441.put(0, t);
    endrule
    rule rule_7524;
        ChannelMessage t;
        t <- mod_5600.get(106);
        mod_4346.put(1, t);
    endrule
    rule rule_7525;
        ChannelMessage t;
        t <- mod_5275.get(0);
        mod_4469.put(4, t);
    endrule
    rule rule_7526;
        ChannelMessage t;
        t <- mod_5632.get(0);
        mod_5125.put(3, t);
    endrule
    rule rule_7527;
        ChannelMessage t;
        t <- mod_5309.get(79);
        mod_3239.put(0, t);
    endrule
    rule rule_7528;
        ChannelMessage t;
        t <- mod_2747.get(2);
        mod_5469.put(0, t);
    endrule
    rule rule_7529;
        ChannelMessage t;
        t <- mod_4715.get(1);
        mod_5313.put(12, t);
    endrule
    rule rule_7530;
        ChannelMessage t;
        t <- mod_5366.get(0);
        mod_4059.put(2, t);
    endrule
    rule rule_7531;
        ChannelMessage t;
        t <- mod_5634.get(0);
        mod_4674.put(3, t);
    endrule
    rule rule_7532;
        ChannelMessage t;
        t <- mod_943.get(1);
        mod_5572.put(0, t);
    endrule
    rule rule_7533;
        ChannelMessage t;
        t <- mod_5623.get(0);
        mod_2050.put(3, t);
    endrule
    rule rule_7534;
        ChannelMessage t;
        t <- mod_2747.get(1);
        mod_5422.put(0, t);
    endrule
    rule rule_7535;
        ChannelMessage t;
        t <- mod_5585.get(0);
        mod_3075.put(3, t);
    endrule
    rule rule_7536;
        ChannelMessage t;
        t <- mod_5467.get(0);
        mod_4141.put(3, t);
    endrule
    rule rule_7537;
        ChannelMessage t;
        t <- mod_5554.get(0);
        mod_1066.put(3, t);
    endrule
    rule rule_7538;
        ChannelMessage t;
        t <- mod_5600.get(7);
        mod_287.put(1, t);
    endrule
    rule rule_7539;
        ChannelMessage t;
        t <- mod_410.get(2);
        mod_5604.put(0, t);
    endrule
    rule rule_7540;
        ChannelMessage t;
        t <- mod_5430.get(0);
        mod_3772.put(3, t);
    endrule
    rule rule_7541;
        ChannelMessage t;
        t <- mod_4264.get(0);
        mod_5313.put(23, t);
    endrule
    rule rule_7542;
        ChannelMessage t;
        t <- mod_5577.get(0);
        mod_205.put(2, t);
    endrule
    rule rule_7543;
        ChannelMessage t;
        t <- mod_369.get(1);
        mod_5599.put(0, t);
    endrule
    rule rule_7544;
        ChannelMessage t;
        t <- mod_1312.get(2);
        mod_5393.put(0, t);
    endrule
    rule rule_7545;
        ChannelMessage t;
        t <- mod_5600.get(30);
        mod_1230.put(1, t);
    endrule
    rule rule_7546;
        ChannelMessage t;
        t <- mod_5309.get(2);
        mod_82.put(0, t);
    endrule
    rule rule_7547;
        ChannelMessage t;
        t <- mod_5309.get(23);
        mod_943.put(0, t);
    endrule
    rule rule_7548;
        ChannelMessage t;
        t <- mod_5488.get(0);
        mod_533.put(3, t);
    endrule
    rule rule_7549;
        ChannelMessage t;
        t <- mod_451.get(2);
        mod_5550.put(0, t);
    endrule
    rule rule_7550;
        ChannelMessage t;
        t <- mod_5279.get(0);
        mod_3772.put(4, t);
    endrule
    rule rule_7551;
        ChannelMessage t;
        t <- mod_5517.get(0);
        mod_574.put(2, t);
    endrule
    rule rule_7552;
        ChannelMessage t;
        t <- mod_5479.get(0);
        mod_615.put(2, t);
    endrule
    rule rule_7553;
        ChannelMessage t;
        t <- mod_3731.get(3);
        mod_5313.put(36, t);
    endrule
    rule rule_7554;
        ChannelMessage t;
        t <- mod_5367.get(0);
        mod_1435.put(4, t);
    endrule
    rule rule_7555;
        ChannelMessage t;
        t <- mod_5600.get(113);
        mod_4633.put(1, t);
    endrule
    rule rule_7556;
        ChannelMessage t;
        t <- mod_3403.get(0);
        mod_5553.put(0, t);
    endrule
    rule rule_7557;
        ChannelMessage t;
        t <- mod_5541.get(0);
        mod_2501.put(3, t);
    endrule
    rule rule_7558;
        ChannelMessage t;
        t <- mod_2214.get(1);
        mod_5313.put(73, t);
    endrule
    rule rule_7559;
        ChannelMessage t;
        t <- mod_4797.get(1);
        mod_5396.put(0, t);
    endrule
    rule rule_7560;
        ChannelMessage t;
        t <- mod_2050.get(0);
        mod_5623.put(0, t);
    endrule
    rule rule_7561;
        ChannelMessage t;
        t <- mod_656.get(1);
        mod_5347.put(0, t);
    endrule
    rule rule_7562;
        ChannelMessage t;
        t <- mod_1558.get(3);
        mod_5589.put(0, t);
    endrule
    rule rule_7563;
        ChannelMessage t;
        t <- mod_5392.get(0);
        mod_287.put(2, t);
    endrule
    rule rule_7564;
        ChannelMessage t;
        t <- mod_5476.get(0);
        mod_3936.put(2, t);
    endrule
    rule rule_7565;
        ChannelMessage t;
        t <- mod_5612.get(0);
        mod_3772.put(2, t);
    endrule
    rule rule_7566;
        ChannelMessage t;
        t <- mod_2091.get(0);
        mod_5569.put(0, t);
    endrule
    rule rule_7567;
        ChannelMessage t;
        t <- mod_5600.get(38);
        mod_1558.put(1, t);
    endrule
    rule rule_7568;
        ChannelMessage t;
        t <- mod_1148.get(0);
        mod_5260.put(0, t);
    endrule
    rule rule_7569;
        ChannelMessage t;
        t <- mod_1517.get(1);
        mod_5314.put(0, t);
    endrule
    rule rule_7570;
        ChannelMessage t;
        t <- mod_5483.get(0);
        mod_697.put(4, t);
    endrule
    rule rule_7571;
        ChannelMessage t;
        t <- mod_5262.get(0);
        mod_1066.put(2, t);
    endrule
    rule rule_7572;
        ChannelMessage t;
        t <- mod_1189.get(0);
        mod_5387.put(0, t);
    endrule
    rule rule_7573;
        ChannelMessage t;
        t <- mod_2255.get(1);
        mod_5364.put(0, t);
    endrule
    rule rule_7574;
        ChannelMessage t;
        t <- mod_5309.get(67);
        mod_2747.put(0, t);
    endrule
    rule rule_7575;
        ChannelMessage t;
        t <- mod_287.get(1);
        mod_5392.put(0, t);
    endrule
    rule rule_7576;
        ChannelMessage t;
        t <- mod_5600.get(23);
        mod_943.put(1, t);
    endrule
    rule rule_7577;
        ChannelMessage t;
        t <- mod_3649.get(3);
        mod_5521.put(0, t);
    endrule
    rule rule_7578;
        ChannelMessage t;
        t <- mod_4920.get(1);
        mod_5276.put(0, t);
    endrule
    rule rule_7579;
        ChannelMessage t;
        t <- mod_5309.get(65);
        mod_2665.put(0, t);
    endrule
    rule rule_7580;
        ChannelMessage t;
        t <- mod_5309.get(84);
        mod_3444.put(0, t);
    endrule
    rule rule_7581;
        ChannelMessage t;
        t <- mod_5472.get(0);
        mod_164.put(2, t);
    endrule
    rule rule_7582;
        ChannelMessage t;
        t <- mod_5309.get(19);
        mod_779.put(0, t);
    endrule
    rule rule_7583;
        ChannelMessage t;
        t <- mod_5346.get(0);
        mod_3608.put(2, t);
    endrule
    rule rule_7584;
        ChannelMessage t;
        t <- mod_5417.get(0);
        mod_1435.put(2, t);
    endrule
    rule rule_7585;
        ChannelMessage t;
        t <- mod_5536.get(0);
        mod_4920.put(3, t);
    endrule
    rule rule_7586;
        ChannelMessage t;
        t <- mod_1189.get(1);
        mod_5313.put(98, t);
    endrule
    rule rule_7587;
        ChannelMessage t;
        t <- mod_5272.get(0);
        mod_82.put(3, t);
    endrule
    rule rule_7588;
        ChannelMessage t;
        t <- mod_2296.get(1);
        mod_5371.put(0, t);
    endrule
    rule rule_7589;
        ChannelMessage t;
        t <- mod_5309.get(114);
        mod_4674.put(0, t);
    endrule
    rule rule_7590;
        ChannelMessage t;
        t <- mod_1353.get(2);
        mod_5513.put(0, t);
    endrule
    rule rule_7591;
        ChannelMessage t;
        t <- mod_1722.get(2);
        mod_5313.put(85, t);
    endrule
    rule rule_7592;
        ChannelMessage t;
        t <- mod_5356.get(0);
        mod_2009.put(2, t);
    endrule
    rule rule_7593;
        ChannelMessage t;
        t <- mod_5043.get(2);
        mod_5253.put(0, t);
    endrule
    rule rule_7594;
        ChannelMessage t;
        t <- mod_5453.get(0);
        mod_2091.put(4, t);
    endrule
    rule rule_7595;
        ChannelMessage t;
        t <- mod_3034.get(0);
        mod_5313.put(53, t);
    endrule
    rule rule_7596;
        ChannelMessage t;
        t <- mod_5309.get(0);
        mod_0.put(0, t);
    endrule
    rule rule_7597;
        ChannelMessage t;
        t <- mod_5495.get(0);
        mod_5255.put(0, t);
    endrule
    rule rule_7598;
        ChannelMessage t;
        t <- mod_5559.get(0);
        mod_4551.put(4, t);
    endrule
    rule rule_7599;
        ChannelMessage t;
        t <- mod_3280.get(2);
        mod_5586.put(0, t);
    endrule
    rule rule_7600;
        ChannelMessage t;
        t <- mod_5443.get(0);
        mod_1189.put(2, t);
    endrule
    rule rule_7601;
        ChannelMessage t;
        t <- mod_5362.get(0);
        mod_738.put(3, t);
    endrule
    rule rule_7602;
        ChannelMessage t;
        t <- mod_5400.get(0);
        mod_3485.put(3, t);
    endrule
    rule rule_7603;
        ChannelMessage t;
        t <- mod_1394.get(2);
        mod_5579.put(0, t);
    endrule
    rule rule_7604;
        ChannelMessage t;
        t <- mod_5248.get(0);
        mod_5580.put(0, t);
    endrule
    rule rule_7605;
        ChannelMessage t;
        t <- mod_5259.get(0);
        mod_3895.put(2, t);
    endrule
    rule rule_7606;
        ChannelMessage t;
        t <- mod_5369.get(0);
        mod_2501.put(2, t);
    endrule
    rule rule_7607;
        ChannelMessage t;
        t <- mod_5600.get(70);
        mod_2870.put(1, t);
    endrule
    rule rule_7608;
        ChannelMessage t;
        t <- mod_5319.get(0);
        mod_3813.put(2, t);
    endrule
    rule rule_7609;
        ChannelMessage t;
        t <- mod_5600.get(111);
        mod_4551.put(1, t);
    endrule
    rule rule_7610;
        ChannelMessage t;
        t <- mod_0.get(2);
        mod_5528.put(0, t);
    endrule
    rule rule_7611;
        ChannelMessage t;
        t <- mod_5478.get(0);
        mod_3977.put(3, t);
    endrule
    rule rule_7612;
        ChannelMessage t;
        t <- mod_5616.get(0);
        mod_4756.put(4, t);
    endrule
    rule rule_7613;
        ChannelMessage t;
        t <- mod_5557.get(0);
        mod_533.put(2, t);
    endrule
    rule rule_7614;
        ChannelMessage t;
        t <- mod_5600.get(42);
        mod_1722.put(1, t);
    endrule
    rule rule_7615;
        ChannelMessage t;
        t <- mod_2214.get(0);
        mod_5416.put(0, t);
    endrule
    rule rule_7616;
        ChannelMessage t;
        t <- mod_5309.get(111);
        mod_4551.put(0, t);
    endrule
    rule rule_7617;
        ChannelMessage t;
        t <- mod_3116.get(2);
        mod_5313.put(51, t);
    endrule
    rule rule_7618;
        ChannelMessage t;
        t <- mod_3198.get(2);
        mod_5313.put(49, t);
    endrule
    rule rule_7619;
        ChannelMessage t;
        t <- mod_123.get(3);
        mod_5500.put(0, t);
    endrule
    rule rule_7620;
        ChannelMessage t;
        t <- mod_41.get(1);
        mod_5431.put(0, t);
    endrule
    rule rule_7621;
        ChannelMessage t;
        t <- mod_5548.get(0);
        mod_328.put(3, t);
    endrule
    rule rule_7622;
        ChannelMessage t;
        t <- mod_5309.get(90);
        mod_3690.put(0, t);
    endrule
    rule rule_7623;
        ChannelMessage t;
        t <- mod_287.get(0);
        mod_5313.put(120, t);
    endrule
    rule rule_7624;
        ChannelMessage t;
        t <- mod_5600.get(62);
        mod_2542.put(1, t);
    endrule
    rule rule_7625;
        ChannelMessage t;
        t <- mod_3649.get(2);
        mod_5313.put(38, t);
    endrule
    rule rule_7626;
        ChannelMessage t;
        t <- mod_656.get(2);
        mod_5370.put(0, t);
    endrule
    rule rule_7627;
        ChannelMessage t;
        t <- mod_4469.get(1);
        mod_5376.put(0, t);
    endrule
    rule rule_7628;
        ChannelMessage t;
        t <- mod_2378.get(3);
        mod_5330.put(0, t);
    endrule
    rule rule_7629;
        ChannelMessage t;
        t <- mod_5600.get(54);
        mod_2214.put(1, t);
    endrule
    rule rule_7630;
        ChannelMessage t;
        t <- mod_5354.get(0);
        mod_4797.put(4, t);
    endrule
    rule rule_7631;
        ChannelMessage t;
        t <- mod_5335.get(0);
        mod_984.put(2, t);
    endrule
    rule rule_7632;
        ChannelMessage t;
        t <- mod_5315.get(0);
        mod_3567.put(4, t);
    endrule
    rule rule_7633;
        ChannelMessage t;
        t <- mod_5309.get(53);
        mod_2173.put(0, t);
    endrule
    rule rule_7634;
        ChannelMessage t;
        t <- mod_3854.get(3);
        mod_5313.put(33, t);
    endrule
    rule rule_7635;
        ChannelMessage t;
        t <- mod_5600.get(51);
        mod_2091.put(1, t);
    endrule
    rule rule_7636;
        ChannelMessage t;
        t <- mod_5603.get(0);
        mod_3526.put(4, t);
    endrule
    rule rule_7637;
        ChannelMessage t;
        t <- mod_5452.get(0);
        mod_369.put(3, t);
    endrule
    rule rule_7638;
        ChannelMessage t;
        t <- mod_5309.get(104);
        mod_4264.put(0, t);
    endrule
    rule rule_7639;
        ChannelMessage t;
        t <- mod_5297.get(0);
        mod_2706.put(2, t);
    endrule
    rule rule_7640;
        ChannelMessage t;
        t <- mod_5600.get(58);
        mod_2378.put(1, t);
    endrule
    rule rule_7641;
        ChannelMessage t;
        t <- mod_4879.get(3);
        mod_5524.put(0, t);
    endrule
    rule rule_7642;
        ChannelMessage t;
        t <- mod_5600.get(41);
        mod_1681.put(1, t);
    endrule
    rule rule_7643;
        ChannelMessage t;
        t <- mod_1435.get(2);
        mod_5283.put(0, t);
    endrule
    rule rule_7644;
        ChannelMessage t;
        t <- mod_5309.get(14);
        mod_574.put(0, t);
    endrule
    rule rule_7645;
        ChannelMessage t;
        t <- mod_1189.get(2);
        mod_5583.put(0, t);
    endrule
    rule rule_7646;
        ChannelMessage t;
        t <- mod_5645.get(0);
        mod_2788.put(2, t);
    endrule
    rule rule_7647;
        ChannelMessage t;
        t <- mod_5309.get(61);
        mod_2501.put(0, t);
    endrule
    rule rule_7648;
        ChannelMessage t;
        t <- mod_5630.get(0);
        mod_1599.put(3, t);
    endrule
    rule rule_7649;
        ChannelMessage t;
        t <- mod_5628.get(0);
        mod_1804.put(4, t);
    endrule
    rule rule_7650;
        ChannelMessage t;
        t <- mod_2214.get(2);
        mod_5590.put(0, t);
    endrule
    rule rule_7651;
        ChannelMessage t;
        t <- mod_5534.get(0);
        mod_3239.put(2, t);
    endrule
    rule rule_7652;
        ChannelMessage t;
        t <- mod_1763.get(1);
        mod_5313.put(84, t);
    endrule
    rule rule_7653;
        ChannelMessage t;
        t <- mod_0.get(0);
        mod_5313.put(127, t);
    endrule
    rule rule_7654;
        ChannelMessage t;
        t <- mod_5600.get(98);
        mod_4018.put(1, t);
    endrule
    rule rule_7655;
        ChannelMessage t;
        t <- mod_5309.get(69);
        mod_2829.put(0, t);
    endrule
    rule rule_7656;
        ChannelMessage t;
        t <- mod_5309.get(95);
        mod_3895.put(0, t);
    endrule
    rule rule_7657;
        ChannelMessage t;
        t <- mod_2665.get(1);
        mod_5313.put(62, t);
    endrule
    rule rule_7658;
        ChannelMessage t;
        t <- mod_5471.get(0);
        mod_1353.put(4, t);
    endrule
    rule rule_7659;
        ChannelMessage t;
        t <- mod_5309.get(127);
        mod_5207.put(0, t);
    endrule
    rule rule_7660;
        ChannelMessage t;
        t <- mod_4387.get(3);
        mod_5512.put(0, t);
    endrule
    rule rule_7661;
        ChannelMessage t;
        t <- mod_2706.get(3);
        mod_5406.put(0, t);
    endrule
    rule rule_7662;
        ChannelMessage t;
        t <- mod_4510.get(2);
        mod_5509.put(0, t);
    endrule
    rule rule_7663;
        ChannelMessage t;
        t <- mod_5600.get(120);
        mod_4920.put(1, t);
    endrule
    rule rule_7664;
        ChannelMessage t;
        t <- mod_5547.get(0);
        mod_902.put(4, t);
    endrule
    rule rule_7665;
        ChannelMessage t;
        t <- mod_1640.get(0);
        mod_5313.put(87, t);
    endrule
    rule rule_7666;
        ChannelMessage t;
        t <- mod_5540.get(0);
        mod_2542.put(4, t);
    endrule
    rule rule_7667;
        ChannelMessage t;
        t <- mod_5558.get(0);
        mod_4510.put(3, t);
    endrule
    rule rule_7668;
        ChannelMessage t;
        t <- mod_5524.get(0);
        mod_4879.put(2, t);
    endrule
    rule rule_7669;
        ChannelMessage t;
        t <- mod_5264.get(0);
        mod_4346.put(2, t);
    endrule
    rule rule_7670;
        ChannelMessage t;
        t <- mod_5462.get(0);
        mod_2378.put(3, t);
    endrule
    rule rule_7671;
        ChannelMessage t;
        t <- mod_5340.get(0);
        mod_3526.put(3, t);
    endrule
    rule rule_7672;
        ChannelMessage t;
        t <- mod_5600.get(75);
        mod_3075.put(1, t);
    endrule
    rule rule_7673;
        ChannelMessage t;
        t <- mod_5491.get(0);
        mod_3649.put(3, t);
    endrule
    rule rule_7674;
        ChannelMessage t;
        t <- mod_5600.get(109);
        mod_4469.put(1, t);
    endrule
    rule rule_7675;
        ChannelMessage t;
        t <- mod_5475.get(0);
        mod_5207.put(3, t);
    endrule
    rule rule_7676;
        ChannelMessage t;
        t <- mod_1189.get(3);
        mod_5443.put(0, t);
    endrule
    rule rule_7677;
        ChannelMessage t;
        t <- mod_4551.get(0);
        mod_5531.put(0, t);
    endrule
    rule rule_7678;
        ChannelMessage t;
        t <- mod_5309.get(123);
        mod_5043.put(0, t);
    endrule
    rule rule_7679;
        ChannelMessage t;
        t <- mod_164.get(3);
        mod_5472.put(0, t);
    endrule
    rule rule_7680;
        ChannelMessage t;
        t <- mod_3075.get(1);
        mod_5466.put(0, t);
    endrule
    rule rule_7681;
        ChannelMessage t;
        t <- mod_164.get(0);
        mod_5489.put(0, t);
    endrule
    rule rule_7682;
        ChannelMessage t;
        t <- mod_779.get(0);
        mod_5639.put(0, t);
    endrule
    rule rule_7683;
        ChannelMessage t;
        t <- mod_1599.get(3);
        mod_5630.put(0, t);
    endrule
    rule rule_7684;
        ChannelMessage t;
        t <- mod_5309.get(124);
        mod_5084.put(0, t);
    endrule
    rule rule_7685;
        ChannelMessage t;
        t <- mod_1476.get(3);
        mod_5313.put(91, t);
    endrule
    rule rule_7686;
        ChannelMessage t;
        t <- mod_2624.get(3);
        mod_5575.put(0, t);
    endrule
    rule rule_7687;
        ChannelMessage t;
        t <- mod_2009.get(0);
        mod_5306.put(0, t);
    endrule
    rule rule_7688;
        ChannelMessage t;
        t <- mod_2829.get(2);
        mod_5591.put(0, t);
    endrule
    rule rule_7689;
        ChannelMessage t;
        t <- mod_5309.get(66);
        mod_2706.put(0, t);
    endrule
    rule rule_7690;
        ChannelMessage t;
        t <- mod_5309.get(126);
        mod_5166.put(0, t);
    endrule
    rule rule_7691;
        ChannelMessage t;
        t <- mod_5448.get(0);
        mod_3198.put(2, t);
    endrule
    rule rule_7692;
        ChannelMessage t;
        t <- mod_5553.get(0);
        mod_3403.put(4, t);
    endrule
    rule rule_7693;
        ChannelMessage t;
        t <- mod_5564.get(0);
        mod_4961.put(2, t);
    endrule
    rule rule_7694;
        ChannelMessage t;
        t <- mod_4428.get(2);
        mod_5250.put(0, t);
    endrule
    rule rule_7695;
        ChannelMessage t;
        t <- mod_1722.get(1);
        mod_5587.put(0, t);
    endrule
    rule rule_7696;
        ChannelMessage t;
        t <- mod_5401.get(0);
        mod_3608.put(4, t);
    endrule
    rule rule_7697;
        ChannelMessage t;
        t <- mod_5635.get(0);
        mod_1558.put(4, t);
    endrule
    rule rule_7698;
        ChannelMessage t;
        t <- mod_2009.get(3);
        mod_5356.put(0, t);
    endrule
    rule rule_7699;
        ChannelMessage t;
        t <- mod_5309.get(13);
        mod_533.put(0, t);
    endrule
    rule rule_7700;
        ChannelMessage t;
        t <- mod_1230.get(2);
        mod_5530.put(0, t);
    endrule
    rule rule_7701;
        ChannelMessage t;
        t <- mod_5600.get(90);
        mod_3690.put(1, t);
    endrule
    rule rule_7702;
        ChannelMessage t;
        t <- mod_2542.get(0);
        mod_5429.put(0, t);
    endrule
    rule rule_7703;
        ChannelMessage t;
        t <- mod_4879.get(0);
        mod_5613.put(0, t);
    endrule
    rule rule_7704;
        ChannelMessage t;
        t <- mod_3485.get(0);
        mod_5588.put(0, t);
    endrule
    rule rule_7705;
        ChannelMessage t;
        t <- mod_5309.get(117);
        mod_4797.put(0, t);
    endrule
    rule rule_7706;
        ChannelMessage t;
        t <- mod_5640.get(0);
        mod_5166.put(3, t);
    endrule
    rule rule_7707;
        ChannelMessage t;
        t <- mod_4920.get(2);
        mod_5294.put(0, t);
    endrule
    rule rule_7708;
        ChannelMessage t;
        t <- mod_1722.get(3);
        mod_5450.put(0, t);
    endrule
    rule rule_7709;
        ChannelMessage t;
        t <- mod_5405.get(0);
        mod_820.put(3, t);
    endrule
    rule rule_7710;
        ChannelMessage t;
        t <- mod_1066.get(0);
        mod_5313.put(101, t);
    endrule
    rule rule_7711;
        ChannelMessage t;
        t <- mod_5600.get(93);
        mod_3813.put(1, t);
    endrule
    rule rule_7712;
        ChannelMessage t;
        t <- mod_5387.get(0);
        mod_1189.put(3, t);
    endrule
    rule rule_7713;
        ChannelMessage t;
        t <- mod_5445.get(0);
        mod_82.put(2, t);
    endrule
    rule rule_7714;
        ChannelMessage t;
        t <- mod_1476.get(1);
        mod_5617.put(0, t);
    endrule
    rule rule_7715;
        ChannelMessage t;
        t <- mod_5600.get(115);
        mod_4715.put(1, t);
    endrule
    rule rule_7716;
        ChannelMessage t;
        t <- mod_5337.get(0);
        mod_246.put(2, t);
    endrule
    rule rule_7717;
        ChannelMessage t;
        t <- mod_5600.get(20);
        mod_820.put(1, t);
    endrule
    rule rule_7718;
        ChannelMessage t;
        t <- mod_5514.get(0);
        mod_2952.put(4, t);
    endrule
    rule rule_7719;
        ChannelMessage t;
        t <- mod_5309.get(52);
        mod_2132.put(0, t);
    endrule
    rule rule_7720;
        ChannelMessage t;
        t <- mod_4059.get(2);
        mod_5366.put(0, t);
    endrule
    rule rule_7721;
        ChannelMessage t;
        t <- mod_5525.get(0);
        mod_4387.put(4, t);
    endrule
    rule rule_7722;
        ChannelMessage t;
        t <- mod_5385.get(0);
        mod_574.put(4, t);
    endrule
    rule rule_7723;
        ChannelMessage t;
        t <- mod_5600.get(99);
        mod_4059.put(1, t);
    endrule
    rule rule_7724;
        ChannelMessage t;
        t <- mod_1886.get(0);
        mod_5602.put(0, t);
    endrule
    rule rule_7725;
        ChannelMessage t;
        t <- mod_5429.get(0);
        mod_2542.put(2, t);
    endrule
    rule rule_7726;
        ChannelMessage t;
        t <- mod_5309.get(70);
        mod_2870.put(0, t);
    endrule
    rule rule_7727;
        ChannelMessage t;
        t <- mod_5440.get(0);
        mod_1886.put(4, t);
    endrule
    rule rule_7728;
        ChannelMessage t;
        t <- mod_5581.get(0);
        mod_1476.put(4, t);
    endrule
    rule rule_7729;
        ChannelMessage t;
        t <- mod_5309.get(81);
        mod_3321.put(0, t);
    endrule
    rule rule_7730;
        ChannelMessage t;
        t <- mod_2665.get(0);
        mod_5595.put(0, t);
    endrule
    rule rule_7731;
        ChannelMessage t;
        t <- mod_5549.get(0);
        mod_861.put(2, t);
    endrule
    rule rule_7732;
        ChannelMessage t;
        t <- mod_5309.get(82);
        mod_3362.put(0, t);
    endrule
    rule rule_7733;
        ChannelMessage t;
        t <- mod_5600.get(100);
        mod_4100.put(1, t);
    endrule
    rule rule_7734;
        ChannelMessage t;
        t <- mod_820.get(3);
        mod_5313.put(107, t);
    endrule
    rule rule_7735;
        ChannelMessage t;
        t <- mod_5357.get(0);
        mod_4961.put(3, t);
    endrule
    rule rule_7736;
        ChannelMessage t;
        t <- mod_5620.get(0);
        mod_5002.put(4, t);
    endrule
    rule rule_7737;
        ChannelMessage t;
        t <- mod_5600.get(35);
        mod_1435.put(1, t);
    endrule
    rule rule_7738;
        ChannelMessage t;
        t <- mod_5309.get(3);
        mod_123.put(0, t);
    endrule
    rule rule_7739;
        ChannelMessage t;
        t <- mod_5600.get(32);
        mod_1312.put(1, t);
    endrule
    rule rule_7740;
        ChannelMessage t;
        t <- mod_1517.get(3);
        mod_5313.put(90, t);
    endrule
    rule rule_7741;
        ChannelMessage t;
        t <- mod_2952.get(0);
        mod_5378.put(0, t);
    endrule
    rule rule_7742;
        ChannelMessage t;
        t <- mod_4592.get(3);
        mod_5442.put(0, t);
    endrule
    rule rule_7743;
        ChannelMessage t;
        t <- mod_5546.get(0);
        mod_5125.put(2, t);
    endrule
    rule rule_7744;
        ChannelMessage t;
        t <- mod_5600.get(18);
        mod_738.put(1, t);
    endrule
    rule rule_7745;
        ChannelMessage t;
        t <- mod_4346.get(3);
        mod_5313.put(21, t);
    endrule
    rule rule_7746;
        ChannelMessage t;
        t <- mod_5600.get(67);
        mod_2747.put(1, t);
    endrule
    rule rule_7747;
        ChannelMessage t;
        t <- mod_2870.get(3);
        mod_5454.put(0, t);
    endrule
    rule rule_7748;
        ChannelMessage t;
        t <- mod_5518.get(0);
        mod_2911.put(2, t);
    endrule
    rule rule_7749;
        ChannelMessage t;
        t <- mod_5473.get(0);
        mod_451.put(4, t);
    endrule
    rule rule_7750;
        ChannelMessage t;
        t <- mod_3731.get(2);
        mod_5496.put(0, t);
    endrule
    rule rule_7751;
        ChannelMessage t;
        t <- mod_4838.get(3);
        mod_5598.put(0, t);
    endrule
    rule rule_7752;
        ChannelMessage t;
        t <- mod_5447.get(0);
        mod_3362.put(2, t);
    endrule
    rule rule_7753;
        ChannelMessage t;
        t <- mod_4100.get(0);
        mod_5499.put(0, t);
    endrule
    rule rule_7754;
        ChannelMessage t;
        t <- mod_4428.get(0);
        mod_5627.put(0, t);
    endrule
    rule rule_7755;
        ChannelMessage t;
        t <- mod_2132.get(1);
        mod_5291.put(0, t);
    endrule
    rule rule_7756;
        ChannelMessage t;
        t <- mod_3731.get(0);
        mod_5642.put(0, t);
    endrule
    rule rule_7757;
        ChannelMessage t;
        t <- mod_5260.get(0);
        mod_1148.put(3, t);
    endrule
    rule rule_7758;
        ChannelMessage t;
        t <- mod_2091.get(2);
        mod_5313.put(76, t);
    endrule
    rule rule_7759;
        ChannelMessage t;
        t <- mod_3075.get(0);
        mod_5464.put(0, t);
    endrule
    rule rule_7760;
        ChannelMessage t;
        t <- mod_5309.get(60);
        mod_2460.put(0, t);
    endrule
    rule rule_7761;
        ChannelMessage t;
        t <- mod_5323.get(0);
        mod_3362.put(3, t);
    endrule
    rule rule_7762;
        ChannelMessage t;
        t <- mod_902.get(3);
        mod_5547.put(0, t);
    endrule
    rule rule_7763;
        ChannelMessage t;
        t <- mod_5263.get(0);
        mod_4387.put(3, t);
    endrule
    rule rule_7764;
        ChannelMessage t;
        t <- mod_1681.get(2);
        mod_5313.put(86, t);
    endrule
    rule rule_7765;
        ChannelMessage t;
        t <- mod_5309.get(39);
        mod_1599.put(0, t);
    endrule
    rule rule_7766;
        ChannelMessage t;
        t <- mod_5309.get(46);
        mod_1886.put(0, t);
    endrule
    rule rule_7767;
        ChannelMessage t;
        t <- mod_5336.get(0);
        mod_4264.put(4, t);
    endrule
    rule rule_7768;
        ChannelMessage t;
        t <- mod_5125.get(2);
        mod_5546.put(0, t);
    endrule
    rule rule_7769;
        ChannelMessage t;
        t <- mod_5420.get(0);
        mod_2214.put(4, t);
    endrule
    rule rule_7770;
        ChannelMessage t;
        t <- mod_861.get(3);
        mod_5549.put(0, t);
    endrule
    rule rule_7771;
        ChannelMessage t;
        t <- mod_5309.get(76);
        mod_3116.put(0, t);
    endrule
    rule rule_7772;
        ChannelMessage t;
        t <- mod_5468.get(0);
        mod_4100.put(4, t);
    endrule
    rule rule_7773;
        ChannelMessage t;
        t <- mod_5578.get(0);
        mod_1599.put(2, t);
    endrule
    rule rule_7774;
        ChannelMessage t;
        t <- mod_5322.get(0);
        mod_3854.put(4, t);
    endrule
    rule rule_7775;
        ChannelMessage t;
        t <- mod_5502.get(0);
        mod_2337.put(2, t);
    endrule
    rule rule_7776;
        ChannelMessage t;
        t <- mod_4059.get(3);
        mod_5560.put(0, t);
    endrule
    rule rule_7777;
        ChannelMessage t;
        t <- mod_943.get(3);
        mod_5313.put(104, t);
    endrule
    rule rule_7778;
        ChannelMessage t;
        t <- mod_123.get(1);
        mod_5313.put(124, t);
    endrule
    rule rule_7779;
        ChannelMessage t;
        t <- mod_3198.get(3);
        mod_5507.put(0, t);
    endrule
    rule rule_7780;
        ChannelMessage t;
        t <- mod_5284.get(0);
        mod_1353.put(3, t);
    endrule
    rule rule_7781;
        ChannelMessage t;
        t <- mod_5509.get(0);
        mod_4510.put(2, t);
    endrule
    rule rule_7782;
        ChannelMessage t;
        t <- mod_4100.get(2);
        mod_5468.put(0, t);
    endrule
    rule rule_7783;
        ChannelMessage t;
        t <- mod_3854.get(1);
        mod_5593.put(0, t);
    endrule
    rule rule_7784;
        ChannelMessage t;
        t <- mod_5301.get(0);
        mod_1271.put(4, t);
    endrule
    rule rule_7785;
        ChannelMessage t;
        t <- mod_5600.get(55);
        mod_2255.put(1, t);
    endrule
    rule rule_7786;
        ChannelMessage t;
        t <- mod_5600.get(91);
        mod_3731.put(1, t);
    endrule
    rule rule_7787;
        ChannelMessage t;
        t <- mod_574.get(2);
        mod_5455.put(0, t);
    endrule
    rule rule_7788;
        ChannelMessage t;
        t <- mod_3895.get(3);
        mod_5544.put(0, t);
    endrule
    rule rule_7789;
        ChannelMessage t;
        t <- mod_5306.get(0);
        mod_2009.put(3, t);
    endrule
    rule rule_7790;
        ChannelMessage t;
        t <- mod_5327.get(0);
        mod_4182.put(3, t);
    endrule
    rule rule_7791;
        ChannelMessage t;
        t <- mod_2788.get(0);
        mod_5645.put(0, t);
    endrule
    rule rule_7792;
        ChannelMessage t;
        t <- mod_5643.get(0);
        mod_4223.put(4, t);
    endrule
    rule rule_7793;
        ChannelMessage t;
        t <- mod_5464.get(0);
        mod_3075.put(2, t);
    endrule
    rule rule_7794;
        ChannelMessage t;
        t <- mod_5470.get(0);
        mod_3116.put(4, t);
    endrule
    rule rule_7795;
        ChannelMessage t;
        t <- mod_5422.get(0);
        mod_2747.put(2, t);
    endrule
    rule rule_7796;
        ChannelMessage t;
        t <- mod_5444.get(0);
        mod_2419.put(2, t);
    endrule
    rule rule_7797;
        ChannelMessage t;
        t <- mod_5310.get(0);
        mod_1927.put(4, t);
    endrule
    rule rule_7798;
        ChannelMessage t;
        t <- mod_2460.get(1);
        mod_5313.put(67, t);
    endrule
    rule rule_7799;
        ChannelMessage t;
        t <- mod_41.get(3);
        mod_5570.put(0, t);
    endrule
    rule rule_7800;
        ChannelMessage t;
        t <- mod_5287.get(0);
        mod_2829.put(2, t);
    endrule
    rule rule_7801;
        ChannelMessage t;
        t <- mod_5309.get(41);
        mod_1681.put(0, t);
    endrule
    rule rule_7802;
        ChannelMessage t;
        t <- mod_5600.get(101);
        mod_4141.put(1, t);
    endrule
    rule rule_7803;
        ChannelMessage t;
        t <- mod_5283.get(0);
        mod_1435.put(3, t);
    endrule
    rule rule_7804;
        ChannelMessage t;
        t <- mod_5304.get(0);
        mod_1312.put(2, t);
    endrule
    rule rule_7805;
        ChannelMessage t;
        t <- mod_5274.get(0);
        mod_5043.put(4, t);
    endrule
    rule rule_7806;
        ChannelMessage t;
        t <- mod_5413.get(0);
        mod_4305.put(2, t);
    endrule
    rule rule_7807;
        ChannelMessage t;
        t <- mod_533.get(1);
        mod_5316.put(0, t);
    endrule
    rule rule_7808;
        ChannelMessage t;
        t <- mod_2460.get(2);
        mod_5338.put(0, t);
    endrule
    rule rule_7809;
        ChannelMessage t;
        t <- mod_4633.get(3);
        mod_5532.put(0, t);
    endrule
    rule rule_7810;
        ChannelMessage t;
        t <- mod_5002.get(2);
        mod_5620.put(0, t);
    endrule
    rule rule_7811;
        ChannelMessage t;
        t <- mod_2542.get(1);
        mod_5286.put(0, t);
    endrule
    rule rule_7812;
        ChannelMessage t;
        t <- mod_3444.get(0);
        mod_5384.put(0, t);
    endrule
    rule rule_7813;
        ChannelMessage t;
        t <- mod_5280.get(0);
        mod_3936.put(3, t);
    endrule
    rule rule_7814;
        ChannelMessage t;
        t <- mod_5551.get(0);
        mod_2296.put(4, t);
    endrule
    rule rule_7815;
        ChannelMessage t;
        t <- mod_5600.get(1);
        mod_41.put(1, t);
    endrule
    rule rule_7816;
        ChannelMessage t;
        t <- mod_5531.get(0);
        mod_4551.put(3, t);
    endrule
    rule rule_7817;
        ChannelMessage t;
        t <- mod_5600.get(26);
        mod_1066.put(1, t);
    endrule
    rule rule_7818;
        ChannelMessage t;
        t <- mod_5609.get(0);
        mod_4182.put(2, t);
    endrule
    rule rule_7819;
        ChannelMessage t;
        t <- mod_738.get(0);
        mod_5381.put(0, t);
    endrule
    rule rule_7820;
        ChannelMessage t;
        t <- mod_1558.get(0);
        mod_5635.put(0, t);
    endrule
    rule rule_7821;
        ChannelMessage t;
        t <- mod_2911.get(0);
        mod_5313.put(56, t);
    endrule
    rule rule_7822;
        ChannelMessage t;
        t <- mod_3936.get(1);
        mod_5476.put(0, t);
    endrule
    rule rule_7823;
        ChannelMessage t;
        t <- mod_3239.get(3);
        mod_5342.put(0, t);
    endrule
    rule rule_7824;
        ChannelMessage t;
        t <- mod_5403.get(0);
        mod_2091.put(2, t);
    endrule
    rule rule_7825;
        ChannelMessage t;
        t <- mod_5309.get(113);
        mod_4633.put(0, t);
    endrule
    rule rule_7826;
        ChannelMessage t;
        t <- mod_2747.get(3);
        mod_5485.put(0, t);
    endrule
    rule rule_7827;
        ChannelMessage t;
        t <- mod_5266.get(0);
        mod_3157.put(3, t);
    endrule
    rule rule_7828;
        ChannelMessage t;
        t <- mod_5309.get(99);
        mod_4059.put(0, t);
    endrule
    rule rule_7829;
        ChannelMessage t;
        t <- mod_5309.get(125);
        mod_5125.put(0, t);
    endrule
    rule rule_7830;
        ChannelMessage t;
        t <- mod_5583.get(0);
        mod_1189.put(4, t);
    endrule
    rule rule_7831;
        ChannelMessage t;
        t <- mod_5257.get(0);
        mod_1599.put(4, t);
    endrule
    rule rule_7832;
        ChannelMessage t;
        t <- mod_5277.get(0);
        mod_1804.put(3, t);
    endrule
    rule rule_7833;
        ChannelMessage t;
        t <- mod_1681.get(3);
        mod_5312.put(0, t);
    endrule
    rule rule_7834;
        ChannelMessage t;
        t <- mod_328.get(1);
        mod_5251.put(0, t);
    endrule
    rule rule_7835;
        ChannelMessage t;
        t <- mod_5622.get(0);
        mod_4879.put(4, t);
    endrule
    rule rule_7836;
        ChannelMessage t;
        t <- mod_3977.get(3);
        mod_5493.put(0, t);
    endrule
    rule rule_7837;
        ChannelMessage t;
        t <- mod_5460.get(0);
        mod_5600.put(0, t);
    endrule
    rule rule_7838;
        ChannelMessage t;
        t <- mod_5621.get(0);
        mod_2911.put(3, t);
    endrule
    rule rule_7839;
        ChannelMessage t;
        t <- mod_5309.get(106);
        mod_4346.put(0, t);
    endrule
    rule rule_7840;
        ChannelMessage t;
        t <- mod_5374.get(0);
        mod_2665.put(3, t);
    endrule
    rule rule_7841;
        ChannelMessage t;
        t <- mod_4510.get(1);
        mod_5368.put(0, t);
    endrule
    rule rule_7842;
        ChannelMessage t;
        t <- mod_574.get(1);
        mod_5313.put(113, t);
    endrule
    rule rule_7843;
        ChannelMessage t;
        t <- mod_943.get(2);
        mod_5490.put(0, t);
    endrule
    rule rule_7844;
        ChannelMessage t;
        t <- mod_5600.get(117);
        mod_4797.put(1, t);
    endrule
    rule rule_7845;
        ChannelMessage t;
        t <- mod_697.get(1);
        mod_5298.put(0, t);
    endrule
    rule rule_7846;
        ChannelMessage t;
        t <- mod_1025.get(1);
        mod_5423.put(0, t);
    endrule
    rule rule_7847;
        ChannelMessage t;
        t <- mod_5309.get(87);
        mod_3567.put(0, t);
    endrule
    rule rule_7848;
        ChannelMessage t;
        t <- mod_41.get(2);
        mod_5313.put(126, t);
    endrule
    rule rule_7849;
        ChannelMessage t;
        t <- mod_5342.get(0);
        mod_3239.put(3, t);
    endrule
    rule rule_7850;
        ChannelMessage t;
        t <- mod_5309.get(112);
        mod_4592.put(0, t);
    endrule
    rule rule_7851;
        ChannelMessage t;
        t <- mod_1886.get(1);
        mod_5440.put(0, t);
    endrule
    rule rule_7852;
        ChannelMessage t;
        t <- mod_5600.get(17);
        mod_697.put(1, t);
    endrule
    rule rule_7853;
        ChannelMessage t;
        t <- mod_2624.get(1);
        mod_5313.put(63, t);
    endrule
    rule rule_7854;
        ChannelMessage t;
        t <- mod_5618.get(0);
        mod_3485.put(4, t);
    endrule
    rule rule_7855;
        ChannelMessage t;
        t <- mod_3157.get(3);
        mod_5355.put(0, t);
    endrule
    rule rule_7856;
        ChannelMessage t;
        t <- mod_2911.get(1);
        mod_5621.put(0, t);
    endrule
    rule rule_7857;
        ChannelMessage t;
        t <- mod_5267.get(0);
        mod_410.put(3, t);
    endrule
    rule rule_7858;
        ChannelMessage t;
        t <- mod_5501.get(0);
        mod_3649.put(4, t);
    endrule
    rule rule_7859;
        ChannelMessage t;
        t <- mod_5600.get(107);
        mod_4387.put(1, t);
    endrule
    rule rule_7860;
        ChannelMessage t;
        t <- mod_5590.get(0);
        mod_2214.put(2, t);
    endrule
    rule rule_7861;
        ChannelMessage t;
        t <- mod_3362.get(3);
        mod_5302.put(0, t);
    endrule
    rule rule_7862;
        ChannelMessage t;
        t <- mod_2132.get(3);
        mod_5313.put(75, t);
    endrule
    rule rule_7863;
        ChannelMessage t;
        t <- mod_5588.get(0);
        mod_3485.put(2, t);
    endrule
    rule rule_7864;
        ChannelMessage t;
        t <- mod_4715.get(3);
        mod_5567.put(0, t);
    endrule
    rule rule_7865;
        ChannelMessage t;
        t <- mod_1394.get(3);
        mod_5592.put(0, t);
    endrule
    rule rule_7866;
        ChannelMessage t;
        t <- mod_5398.get(0);
        mod_3567.put(2, t);
    endrule
    rule rule_7867;
        ChannelMessage t;
        t <- mod_5600.get(72);
        mod_2952.put(1, t);
    endrule
    rule rule_7868;
        ChannelMessage t;
        t <- mod_123.get(0);
        mod_5328.put(0, t);
    endrule
    rule rule_7869;
        ChannelMessage t;
        t <- mod_5636.get(0);
        mod_3034.put(4, t);
    endrule
    rule rule_7870;
        ChannelMessage t;
        t <- mod_5600.get(104);
        mod_4264.put(1, t);
    endrule
    rule rule_7871;
        ChannelMessage t;
        t <- mod_1886.get(3);
        mod_5542.put(0, t);
    endrule
    rule rule_7872;
        ChannelMessage t;
        t <- mod_4715.get(0);
        mod_5373.put(0, t);
    endrule
    rule rule_7873;
        ChannelMessage t;
        t <- mod_4674.get(3);
        mod_5375.put(0, t);
    endrule
    rule rule_7874;
        ChannelMessage t;
        t <- mod_5523.get(0);
        mod_5313.put(128, t);
    endrule
    rule rule_7875;
        ChannelMessage t;
        t <- mod_5343.get(0);
        mod_615.put(4, t);
    endrule
    rule rule_7876;
        ChannelMessage t;
        t <- mod_3526.get(2);
        mod_5340.put(0, t);
    endrule
    rule rule_7877;
        ChannelMessage t;
        t <- mod_3034.get(1);
        mod_5252.put(0, t);
    endrule
    rule rule_7878;
        ChannelMessage t;
        t <- mod_5309.get(1);
        mod_41.put(0, t);
    endrule
    rule rule_7879;
        ChannelMessage t;
        t <- mod_5600.get(69);
        mod_2829.put(1, t);
    endrule
    rule rule_7880;
        ChannelMessage t;
        t <- mod_5372.get(1);
        mod_5495.put(0, t);
    endrule
    rule rule_7881;
        ChannelMessage t;
        t <- mod_5573.get(0);
        mod_2173.put(3, t);
    endrule
    rule rule_7882;
        ChannelMessage t;
        t <- mod_4633.get(1);
        mod_5313.put(14, t);
    endrule
    rule rule_7883;
        ChannelMessage t;
        t <- mod_4469.get(2);
        mod_5313.put(18, t);
    endrule
    rule rule_7884;
        ChannelMessage t;
        t <- mod_5289.get(0);
        mod_4018.put(4, t);
    endrule
    rule rule_7885;
        ChannelMessage t;
        t <- mod_5309.get(73);
        mod_2993.put(0, t);
    endrule
    rule rule_7886;
        ChannelMessage t;
        t <- mod_5406.get(0);
        mod_2706.put(4, t);
    endrule
    rule rule_7887;
        ChannelMessage t;
        t <- mod_5597.get(0);
        mod_1148.put(4, t);
    endrule
    rule rule_7888;
        ChannelMessage t;
        t <- mod_5043.get(3);
        mod_5313.put(4, t);
    endrule
    rule rule_7889;
        ChannelMessage t;
        t <- mod_4510.get(0);
        mod_5313.put(17, t);
    endrule
    rule rule_7890;
        ChannelMessage t;
        t <- mod_3157.get(0);
        mod_5647.put(0, t);
    endrule
    rule rule_7891;
        ChannelMessage t;
        t <- mod_5207.get(0);
        mod_5313.put(0, t);
    endrule
    rule rule_7892;
        ChannelMessage t;
        t <- mod_5600.get(47);
        mod_1927.put(1, t);
    endrule
    rule rule_7893;
        ChannelMessage t;
        t <- mod_3690.get(0);
        mod_5607.put(0, t);
    endrule
    rule rule_7894;
        ChannelMessage t;
        t <- mod_1025.get(3);
        mod_5313.put(102, t);
    endrule
    rule rule_7895;
        ChannelMessage t;
        t <- mod_5570.get(0);
        mod_41.put(4, t);
    endrule
    rule rule_7896;
        ChannelMessage t;
        t <- mod_5309.get(24);
        mod_984.put(0, t);
    endrule
    rule rule_7897;
        ChannelMessage t;
        t <- mod_1435.get(3);
        mod_5313.put(92, t);
    endrule
    rule rule_7898;
        ChannelMessage t;
        t <- mod_5002.get(1);
        mod_5388.put(0, t);
    endrule
    rule rule_7899;
        ChannelMessage t;
        t <- mod_5309.get(48);
        mod_1968.put(0, t);
    endrule
    rule rule_7900;
        ChannelMessage t;
        t <- mod_5309.get(100);
        mod_4100.put(0, t);
    endrule
    rule rule_7901;
        ChannelMessage t;
        t <- mod_5600.get(81);
        mod_3321.put(1, t);
    endrule
    rule rule_7902;
        ChannelMessage t;
        t <- mod_2706.get(2);
        mod_5297.put(0, t);
    endrule
    rule rule_7903;
        ChannelMessage t;
        t <- mod_4141.get(1);
        mod_5410.put(0, t);
    endrule
    rule rule_7904;
        ChannelMessage t;
        t <- mod_3075.get(3);
        mod_5313.put(52, t);
    endrule
    rule rule_7905;
        ChannelMessage t;
        t <- mod_4674.get(0);
        mod_5634.put(0, t);
    endrule
    rule rule_7906;
        ChannelMessage t;
        t <- mod_3157.get(2);
        mod_5313.put(50, t);
    endrule
    rule rule_7907;
        ChannelMessage t;
        t <- mod_1066.get(2);
        mod_5308.put(0, t);
    endrule
    rule rule_7908;
        ChannelMessage t;
        t <- mod_2870.get(1);
        mod_5629.put(0, t);
    endrule
    rule rule_7909;
        ChannelMessage t;
        t <- mod_1804.get(1);
        mod_5313.put(83, t);
    endrule
    rule rule_7910;
        ChannelMessage t;
        t <- mod_5365.get(0);
        mod_2378.put(4, t);
    endrule
    rule rule_7911;
        ChannelMessage t;
        t <- mod_5397.get(0);
        mod_4838.put(4, t);
    endrule
    rule rule_7912;
        ChannelMessage t;
        t <- mod_5481.get(0);
        mod_5526.put(0, t);
    endrule
    rule rule_7913;
        ChannelMessage t;
        t <- mod_5511.get(0);
        mod_4223.put(3, t);
    endrule
    rule rule_7914;
        ChannelMessage t;
        t <- mod_861.get(1);
        mod_5285.put(0, t);
    endrule
    rule rule_7915;
        ChannelMessage t;
        t <- mod_1353.get(0);
        mod_5284.put(0, t);
    endrule
    rule rule_7916;
        ChannelMessage t;
        t <- mod_3362.get(1);
        mod_5447.put(0, t);
    endrule
    rule rule_7917;
        ChannelMessage t;
        t <- mod_5600.get(97);
        mod_3977.put(1, t);
    endrule
    rule rule_7918;
        ChannelMessage t;
        t <- mod_5600.get(124);
        mod_5084.put(1, t);
    endrule
    rule rule_7919;
        ChannelMessage t;
        t <- mod_3936.get(0);
        mod_5256.put(0, t);
    endrule
    rule rule_7920;
        ChannelMessage t;
        t <- mod_3567.get(2);
        mod_5398.put(0, t);
    endrule
    rule rule_7921;
        ChannelMessage t;
        t <- mod_5312.get(0);
        mod_1681.put(3, t);
    endrule
    rule rule_7922;
        ChannelMessage t;
        t <- mod_3731.get(1);
        mod_5487.put(0, t);
    endrule
    rule rule_7923;
        ChannelMessage t;
        t <- mod_5309.get(50);
        mod_2050.put(0, t);
    endrule
    rule rule_7924;
        ChannelMessage t;
        t <- mod_5317.get(0);
        mod_4715.put(3, t);
    endrule
    rule rule_7925;
        ChannelMessage t;
        t <- mod_5307.get(0);
        mod_738.put(4, t);
    endrule
    rule rule_7926;
        ChannelMessage t;
        t <- mod_5084.get(1);
        mod_5418.put(0, t);
    endrule
    rule rule_7927;
        ChannelMessage t;
        t <- mod_5309.get(78);
        mod_3198.put(0, t);
    endrule
    rule rule_7928;
        ChannelMessage t;
        t <- mod_5309.get(54);
        mod_2214.put(0, t);
    endrule
    rule rule_7929;
        ChannelMessage t;
        t <- mod_5383.get(0);
        mod_3198.put(4, t);
    endrule
    rule rule_7930;
        ChannelMessage t;
        t <- mod_410.get(1);
        mod_5399.put(0, t);
    endrule
    rule rule_7931;
        ChannelMessage t;
        t <- mod_2337.get(2);
        mod_5522.put(0, t);
    endrule
    rule rule_7932;
        ChannelMessage t;
        t <- mod_3772.get(0);
        mod_5279.put(0, t);
    endrule
    rule rule_7933;
        ChannelMessage t;
        t <- mod_5538.get(0);
        mod_1968.put(3, t);
    endrule
    rule rule_7934;
        ChannelMessage t;
        t <- mod_5600.get(15);
        mod_615.put(1, t);
    endrule
    rule rule_7935;
        ChannelMessage t;
        t <- mod_5309.get(15);
        mod_615.put(0, t);
    endrule
    rule rule_7936;
        ChannelMessage t;
        t <- mod_5600.get(57);
        mod_2337.put(1, t);
    endrule
    rule rule_7937;
        ChannelMessage t;
        t <- mod_5598.get(0);
        mod_4838.put(2, t);
    endrule
    rule rule_7938;
        ChannelMessage t;
        t <- mod_1763.get(3);
        mod_5409.put(0, t);
    endrule
    rule rule_7939;
        ChannelMessage t;
        t <- mod_1763.get(2);
        mod_5290.put(0, t);
    endrule
    rule rule_7940;
        ChannelMessage t;
        t <- mod_5552.get(0);
        mod_5002.put(3, t);
    endrule
    rule rule_7941;
        ChannelMessage t;
        t <- mod_615.get(3);
        mod_5474.put(0, t);
    endrule
    rule rule_7942;
        ChannelMessage t;
        t <- mod_5446.get(0);
        mod_5125.put(4, t);
    endrule
    rule rule_7943;
        ChannelMessage t;
        t <- mod_5566.get(0);
        mod_164.put(3, t);
    endrule
    rule rule_7944;
        ChannelMessage t;
        t <- mod_1558.get(2);
        mod_5269.put(0, t);
    endrule
    rule rule_7945;
        ChannelMessage t;
        t <- mod_4756.get(1);
        mod_5278.put(0, t);
    endrule
    rule rule_7946;
        ChannelMessage t;
        t <- mod_5321.get(0);
        mod_2009.put(4, t);
    endrule
    rule rule_7947;
        ChannelMessage t;
        t <- mod_5384.get(0);
        mod_3444.put(4, t);
    endrule
    rule rule_7948;
        ChannelMessage t;
        t <- mod_5399.get(0);
        mod_410.put(4, t);
    endrule
    rule rule_7949;
        ChannelMessage t;
        t <- mod_5412.get(0);
        mod_2993.put(2, t);
    endrule
    rule rule_7950;
        ChannelMessage t;
        t <- mod_779.get(3);
        mod_5313.put(108, t);
    endrule
    rule rule_7951;
        ChannelMessage t;
        t <- mod_2501.get(3);
        mod_5363.put(0, t);
    endrule
    rule rule_7952;
        ChannelMessage t;
        t <- mod_3116.get(3);
        mod_5543.put(0, t);
    endrule

endmodule
endpackage
