// Currently we access the set / frame by using [0000,SetBit,FrameBit] as a single value

package PMU;

import FIFO::*;
import Types::*;
import Vector::*;
import RegFile::*;
import BankedMemory::*;
import Parameters::*;
import SetFreeList::*;
import SetUsageTracker::*;

// Tracking the current storage location
typedef struct {
    SETS_LOG set;
    FRAMES_PER_SET_LOG frame;
    Bool valid;
} StorageLocation deriving(Bits, Eq);

typedef struct {
  Vector#(MAX_ENTRIES, StorageLocation) vec;
  UInt#(TLog#(MAX_ENTRIES)) next_idx;
} TokenMapping deriving (Bits, Eq);

// Interface that just exposes the modules existence
interface PMU_IFC;
endinterface

// PMU module that processes between the FIFOs
module mkPMU#(
    FIFO#(ChannelMessage) data_in,      // Values come in here
    FIFO#(ChannelMessage) token_out,    // Generated tokens go out here
    FIFO#(ChannelMessage) token_in,     // Tokens come back in here
    FIFO#(ChannelMessage) data_out,     // Retrieved values go out here
    Int#(32) rank_in                    // Rank of the current tile
)(PMU_IFC);
    
    // Only internal state needed is the storage FIFO and token counter
    BankedMemory_IFC mem <- mkBankedMemory;
    SetFreeList_IFC free_list <- mkSetFreeList;
    SetUsageTracker_IFC usage_tracker <- mkSetUsageTracker;
    Reg#(StorageLocation) curr_loc <- mkReg(StorageLocation { set: 0, frame: 0, valid: False });
    Reg#(Int#(32)) rank <- mkReg(rank_in);
    Reg#(Scalar) token_counter <- mkReg(0);
    RegFile#(Scalar, TokenMapping) token_table <- mkRegFile(0, fromInteger(valueOf(MAX_ENTRIES) - 1));
    let frame_width = valueOf(TLog#(FRAMES_PER_SET));
    let set_width = valueOf(TLog#(SETS));
    Reg#(Maybe#(Scalar)) load_token <- mkReg(tagged Invalid);
    Reg#(UInt#(TLog#(MAX_ENTRIES))) load_idx <- mkReg(0);
    
    Reg#(Bool) token_table_initialized <- mkReg(False);
    Reg#(Scalar) init_counter <- mkReg(0);
    rule init_token_table (!token_table_initialized);
        TokenMapping tm;
        tm.vec = replicate(StorageLocation { set: 0, frame: 0, valid: False });
        tm.next_idx = 0;
        token_table.upd(init_counter, tm);

        if (init_counter == fromInteger(valueOf(MAX_ENTRIES) - 1)) begin
            token_table_initialized <= True;
        end else begin
            init_counter <= init_counter + 1;
        end
    endrule

    rule store_tile (token_table_initialized);
        let d_in = data_in.first;
        data_in.deq;

        case (d_in) matches
            tagged Tag_Data {.tt, .st}: begin
                case (tt) matches
                    tagged Tag_Tile .tile: begin
                        let new_st = st;
                        let emit_token = False;
                        if (st >= rank) begin
                            new_st = st - rank;
                            emit_token = True;
                        end

                        StorageLocation new_loc = curr_loc;
                        StorageLocation storage_location = curr_loc;

                        if (!curr_loc.valid) begin
                            let mset <- free_list.allocSet();
                            case (mset) matches
                                tagged Valid .set: begin
                                    mem.write(set, 0, TaggedTile { t: tile, st: st });
                                    usage_tracker.setFrame(set, 1);

                                    FRAMES_PER_SET_LOG zero_frame = 0;
                                    storage_location = StorageLocation { set: set, frame: 0, valid: True };
                                    new_loc = StorageLocation { set: set, frame: 1, valid: True };
                                end
                                default: begin
                                    $display("***** Out of memory *****");
                                    $finish;
                                end
                            endcase
                        end else begin
                            let set = curr_loc.set;
                            let frame = curr_loc.frame;
                            storage_location = curr_loc;

                            mem.write(set, frame, TaggedTile { t: tile, st: st });
                            let full <- usage_tracker.incFrame(set);

                            new_loc = StorageLocation {
                                set: set,
                                frame: frame + 1,
                                valid: !full
                            };
                        end

                        let tm = token_table.sub(token_counter);
                        tm.vec[tm.next_idx] = storage_location;
                        tm.next_idx = tm.next_idx + 1;
                        token_table.upd(token_counter, tm);

                        if (emit_token) begin
                            let token_to_emit = token_counter;
                            token_counter <= token_counter + 1;
                            token_out.enq(tagged Tag_Data tuple2(tagged Tag_Scalar token_to_emit, new_st));
                        end
                        curr_loc <= new_loc;
                    end
                    tagged Tag_Ref .r: begin
                        $display("[ERROR]: Reference received in data input");
                        $finish(0);
                    end
                    tagged Tag_Scalar .scalar: begin
                        $display("[ERROR]: Scalar received in data input");
                        $finish(0);
                    end
                endcase
            end
            tagged Tag_Instruction .ip: begin
                $display("[ERROR]: Instruction received in data input"); // TODO: Should be able to accept incoming config
                $finish(0);
            end
            tagged Tag_EndToken .et: begin
                token_out.enq(tagged Tag_EndToken et);
                $display("End token received in store");
            end
        endcase
    endrule

    // Rule to handle token retrievals: find matching value and return it
    rule start_load_tile (load_token == tagged Invalid);
        let token_msg = token_in.first;
        token_in.deq;
        
        case (token_msg) matches
            tagged Tag_Data {.tt, .st}: begin
                case (tt) matches
                    tagged Tag_Scalar .token_input: begin
                        load_token <= tagged Valid token_input;
                        load_idx <= 0;
                    end
                    default: begin
                        $display("[ERROR]: Expected scalar token");
                        $finish(0);
                    end
                endcase
            end
            tagged Tag_EndToken .et: begin
                // Print the state of the memory being used
                for (Integer i = 0; i < valueOf(SETS); i = i + 1) begin
                    // Check if set is valid
                    if (!free_list.isSetFree(fromInteger(i))) begin
                        $display("[MEMORY USAGE]: Set %d: %d frames used", i, usage_tracker.getCount(fromInteger(i)));
                    end else begin
                        $display("[MEMORY USAGE]: Set %d: No frames used", i);
                    end
                end
                data_out.enq(tagged Tag_EndToken et);
                $display("End token received");
            end
            default: begin
                $display("[ERROR]: Expected data message with token");
                $finish(0);
            end
        endcase
    endrule

    rule continue_load_tile (isValid(load_token));
        $display("[DEBUG]: Continuing load tile %d", fromMaybe(0, load_token));
        let tm = token_table.sub(fromMaybe(0, load_token));
        if (load_idx < tm.next_idx) begin
            let loc = tm.vec[load_idx];
            let set = loc.set;
            let frame = loc.frame;
            let tile = mem.read(set, frame);
            data_out.enq(tagged Tag_Data tuple2(tagged Tag_Tile tile.t, tile.st));
            if (load_idx == tm.next_idx - 1) begin
                load_token <= tagged Invalid;
                load_idx <= 0;
            end else begin
                load_idx <= load_idx + 1;
            end
        end
    endrule

endmodule

endpackage