package Step;
import Operation::*;
import Types::*;
import Vector::*;
import FShow::*;
import Debug::*;
import PMU::*;
import RamulatorArbiter::*;
import RandomLoad::*;

(* synthesize *)
module mkHypernode (Operation_IFC);
    Operation_IFC mod_4839_inner <- mkReshape(2, 64);
    Operation_IFC mod_4839 <- mkDebugOperation(mod_4839_inner, "mod_4839");
    Operation_IFC mod_4840_inner <- mkFlatten(1);
    Operation_IFC mod_4840 <- mkDebugOperation(mod_4840_inner, "mod_4840");
    Operation_IFC mod_4841_inner <- mkFlatten(2);
    Operation_IFC mod_4841 <- mkDebugOperation(mod_4841_inner, "mod_4841");
    Operation_IFC mod_4842_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4842 <- mkDebugOperation(mod_4842_inner, "mod_4842");
    Broadcast_IFC#(4) mod_4843_inner <- mkBroadcast(4);
    Operation_IFC mod_4843 <- mkDebugOperation(mod_4843_inner.op, "mod_4843");
    PMU_IFC mod_4844_bufferize <- mkPMU(2);
    Operation_IFC mod_4844_inner = mod_4844_bufferize.operation;
    Operation_IFC mod_4844 <- mkDebugOperation(mod_4844_inner, "mod_4844");
    Broadcast_IFC#(2) mod_4845_inner <- mkBroadcast(2);
    Operation_IFC mod_4845 <- mkDebugOperation(mod_4845_inner.op, "mod_4845");
    PMU_IFC mod_4846_bufferize <- mkPMU(1);
    Operation_IFC mod_4846_inner = mod_4846_bufferize.operation;
    Operation_IFC mod_4846 <- mkDebugOperation(mod_4846_inner, "mod_4846");
    Operation_IFC mod_4847_inner <- mkBinaryMap(1038, matmul_t_tile);
    Operation_IFC mod_4847 <- mkDebugOperation(mod_4847_inner, "mod_4847");
    Operation_IFC mod_4848_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4848 <- mkDebugOperation(mod_4848_inner, "mod_4848");
    Operation_IFC mod_4849_inner <- mkBinaryMap(1806, mul_tile);
    Operation_IFC mod_4849 <- mkDebugOperation(mod_4849_inner, "mod_4849");
    PMU_IFC mod_4850_bufferize <- mkPMU(1);
    Operation_IFC mod_4850_inner = mod_4850_bufferize.operation;
    Operation_IFC mod_4850 <- mkDebugOperation(mod_4850_inner, "mod_4850");
    Operation_IFC mod_4851_inner <- mkBinaryMap(2327, matmul_t_tile);
    Operation_IFC mod_4851 <- mkDebugOperation(mod_4851_inner, "mod_4851");
    Operation_IFC mod_4852_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4852 <- mkDebugOperation(mod_4852_inner, "mod_4852");
    Operation_IFC mod_4853_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_4853 <- mkDebugOperation(mod_4853_inner, "mod_4853");
    Operation_IFC mod_4854_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_4854 <- mkDebugOperation(mod_4854_inner, "mod_4854");
    Operation_IFC mod_4855_inner <- mkBinaryMap(2705, mul_tile);
    Operation_IFC mod_4855 <- mkDebugOperation(mod_4855_inner, "mod_4855");
    PMU_IFC mod_4856_bufferize <- mkPMU(1);
    Operation_IFC mod_4856_inner = mod_4856_bufferize.operation;
    Operation_IFC mod_4856 <- mkDebugOperation(mod_4856_inner, "mod_4856");
    PMU_IFC mod_4857_bufferize <- mkPMU(2);
    Operation_IFC mod_4857_inner = mod_4857_bufferize.operation;
    Operation_IFC mod_4857 <- mkDebugOperation(mod_4857_inner, "mod_4857");
    PMU_IFC mod_4858_bufferize <- mkPMU(2);
    Operation_IFC mod_4858_inner = mod_4858_bufferize.operation;
    Operation_IFC mod_4858 <- mkDebugOperation(mod_4858_inner, "mod_4858");
    Operation_IFC mod_4859_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4859 <- mkDebugOperation(mod_4859_inner, "mod_4859");
    Operation_IFC mod_4860_inner <- mkFlatten(1);
    Operation_IFC mod_4860 <- mkDebugOperation(mod_4860_inner, "mod_4860");
    Operation_IFC mod_4861_inner <- mkFlatten(0);
    Operation_IFC mod_4861 <- mkDebugOperation(mod_4861_inner, "mod_4861");
    Operation_IFC mod_4862_inner <- mkRepeatStatic(3);
    Operation_IFC mod_4862 <- mkDebugOperation(mod_4862_inner, "mod_4862");
    Operation_IFC mod_4863_inner <- mkUnaryMap(1678, silu_tile);
    Operation_IFC mod_4863 <- mkDebugOperation(mod_4863_inner, "mod_4863");
    Operation_IFC mod_4864_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_4864 <- mkDebugOperation(mod_4864_inner, "mod_4864");
    Operation_IFC mod_4865_inner <- mkBinaryMap(1550, matmul_t_tile);
    Operation_IFC mod_4865 <- mkDebugOperation(mod_4865_inner, "mod_4865");
    PMU_IFC mod_4866_bufferize <- mkPMU(2);
    Operation_IFC mod_4866_inner = mod_4866_bufferize.operation;
    Operation_IFC mod_4866 <- mkDebugOperation(mod_4866_inner, "mod_4866");
    Operation_IFC mod_4867_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4867 <- mkDebugOperation(mod_4867_inner, "mod_4867");
    Operation_IFC mod_4868_inner <- mkFlatten(1);
    Operation_IFC mod_4868 <- mkDebugOperation(mod_4868_inner, "mod_4868");
    Operation_IFC mod_4869_inner <- mkFlatten(0);
    Operation_IFC mod_4869 <- mkDebugOperation(mod_4869_inner, "mod_4869");
    PMU_IFC mod_4870_bufferize <- mkPMU(1);
    Operation_IFC mod_4870_inner = mod_4870_bufferize.operation;
    Operation_IFC mod_4870 <- mkDebugOperation(mod_4870_inner, "mod_4870");
    Operation_IFC mod_4871_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4871 <- mkDebugOperation(mod_4871_inner, "mod_4871");
    PMU_IFC mod_4872_bufferize <- mkPMU(2);
    Operation_IFC mod_4872_inner = mod_4872_bufferize.operation;
    Operation_IFC mod_4872 <- mkDebugOperation(mod_4872_inner, "mod_4872");
    Operation_IFC mod_4873_inner <- mkRepeatStatic(8);
    Operation_IFC mod_4873 <- mkDebugOperation(mod_4873_inner, "mod_4873");
    Operation_IFC mod_4874_inner <- mkFlatten(1);
    Operation_IFC mod_4874 <- mkDebugOperation(mod_4874_inner, "mod_4874");
    Operation_IFC mod_4875_inner <- mkFlatten(0);
    Operation_IFC mod_4875 <- mkDebugOperation(mod_4875_inner, "mod_4875");
    Operation_IFC mod_4876_inner <- mkRepeatStatic(16);
    Operation_IFC mod_4876 <- mkDebugOperation(mod_4876_inner, "mod_4876");
    Operation_IFC mod_4877_inner <- mkRepeatStatic(2);
    Operation_IFC mod_4877 <- mkDebugOperation(mod_4877_inner, "mod_4877");
    PMU_IFC mod_4878_bufferize <- mkPMU(2);
    Operation_IFC mod_4878_inner = mod_4878_bufferize.operation;
    Operation_IFC mod_4878 <- mkDebugOperation(mod_4878_inner, "mod_4878");
    rule rule_6255;
        ChannelMessage t;
        t <- mod_4861.get(0);
        mod_4860.put(0, t);
    endrule
    rule rule_6256;
        ChannelMessage t;
        t <- mod_4856.get(1);
        mod_4854.put(1, t);
    endrule
    rule rule_6257;
        ChannelMessage t;
        t <- mod_4849.get(0);
        mod_4850.put(0, t);
    endrule
    rule rule_6258;
        ChannelMessage t;
        t <- mod_4843.get(3);
        mod_4844.put(0, t);
    endrule
    rule rule_6259;
        ChannelMessage t;
        t <- mod_4844.get(1);
        mod_4845.put(0, t);
    endrule
    rule rule_6260;
        ChannelMessage t;
        t <- mod_4859.get(0);
        mod_4858.put(1, t);
    endrule
    rule rule_6261;
        ChannelMessage t;
        t <- mod_4840.get(0);
        mod_4841.put(0, t);
    endrule
    rule rule_6262;
        ChannelMessage t;
        t <- mod_4870.get(0);
        mod_4871.put(0, t);
    endrule
    rule rule_6263;
        ChannelMessage t;
        t <- mod_4873.get(0);
        mod_4872.put(1, t);
    endrule
    rule rule_6264;
        ChannelMessage t;
        t <- mod_4853.get(1);
        mod_4854.put(0, t);
    endrule
    rule rule_6265;
        ChannelMessage t;
        t <- mod_4864.get(0);
        mod_4863.put(0, t);
    endrule
    rule rule_6266;
        ChannelMessage t;
        t <- mod_4853.get(0);
        mod_4857.put(0, t);
    endrule
    rule rule_6267;
        ChannelMessage t;
        t <- mod_4857.get(0);
        mod_4857.put(1, t);
    endrule
    rule rule_6268;
        ChannelMessage t;
        t <- mod_4870.get(1);
        mod_4865.put(0, t);
    endrule
    rule rule_6269;
        ChannelMessage t;
        t <- mod_4871.get(0);
        mod_4870.put(1, t);
    endrule
    rule rule_6270;
        ChannelMessage t;
        t <- mod_4866.get(0);
        mod_4867.put(0, t);
    endrule
    rule rule_6271;
        ChannelMessage t;
        t <- mod_4872.get(0);
        mod_4873.put(0, t);
    endrule
    rule rule_6272;
        ChannelMessage t;
        t <- mod_4850.get(0);
        mod_4862.put(0, t);
    endrule
    rule rule_6273;
        ChannelMessage t;
        t <- mod_4878.get(1);
        mod_4842.put(1, t);
    endrule
    rule rule_6274;
        ChannelMessage t;
        t <- mod_4872.get(1);
        mod_4847.put(1, t);
    endrule
    rule rule_6275;
        ChannelMessage t;
        t <- mod_4875.get(0);
        mod_4874.put(0, t);
    endrule
    rule rule_6276;
        ChannelMessage t;
        t <- mod_4842.get(1);
        mod_4843.put(0, t);
    endrule
    rule rule_6277;
        ChannelMessage t;
        t <- mod_4867.get(0);
        mod_4866.put(1, t);
    endrule
    rule rule_6278;
        ChannelMessage t;
        t <- mod_4878.get(0);
        mod_4878.put(1, t);
    endrule
    rule rule_6279;
        ChannelMessage t;
        t <- mod_4851.get(0);
        mod_4852.put(0, t);
    endrule
    rule rule_6280;
        ChannelMessage t;
        t <- mod_4848.get(0);
        mod_4849.put(0, t);
    endrule
    rule rule_6281;
        ChannelMessage t;
        t <- mod_4850.get(1);
        mod_4851.put(0, t);
    endrule
    rule rule_6282;
        ChannelMessage t;
        t <- mod_4857.get(1);
        mod_4853.put(1, t);
    endrule
    rule rule_6283;
        ChannelMessage t;
        t <- mod_4852.get(0);
        mod_4853.put(0, t);
    endrule
    rule rule_6284;
        ChannelMessage t;
        t <- mod_4842.get(0);
        mod_4878.put(0, t);
    endrule
    rule rule_6285;
        ChannelMessage t;
        t <- mod_4854.get(0);
        mod_4856.put(0, t);
    endrule
    rule rule_6286;
        ChannelMessage t;
        t <- mod_4858.get(1);
        mod_4851.put(1, t);
    endrule
    rule rule_6287;
        ChannelMessage t;
        t <- mod_4868.get(0);
        mod_4866.put(0, t);
    endrule
    rule rule_6288;
        ChannelMessage t;
        t <- mod_4863.get(0);
        mod_4849.put(1, t);
    endrule
    rule rule_6289;
        ChannelMessage t;
        t <- mod_4869.get(0);
        mod_4868.put(0, t);
    endrule
    rule rule_6290;
        ChannelMessage t;
        t <- mod_4839.get(0);
        mod_4840.put(0, t);
    endrule
    rule rule_6291;
        ChannelMessage t;
        t <- mod_4876.get(0);
        mod_4846.put(1, t);
    endrule
    rule rule_6292;
        ChannelMessage t;
        t <- mod_4854.get(1);
        mod_4855.put(1, t);
    endrule
    rule rule_6293;
        ChannelMessage t;
        t <- mod_4874.get(0);
        mod_4872.put(0, t);
    endrule
    rule rule_6294;
        ChannelMessage t;
        t <- mod_4846.get(1);
        mod_4847.put(0, t);
    endrule
    rule rule_6295;
        ChannelMessage t;
        t <- mod_4847.get(0);
        mod_4848.put(0, t);
    endrule
    rule rule_6296;
        ChannelMessage t;
        t <- mod_4860.get(0);
        mod_4858.put(0, t);
    endrule
    rule rule_6297;
        ChannelMessage t;
        t <- mod_4865.get(0);
        mod_4864.put(0, t);
    endrule
    rule rule_6298;
        ChannelMessage t;
        t <- mod_4846.get(0);
        mod_4876.put(0, t);
    endrule
    rule rule_6299;
        ChannelMessage t;
        t <- mod_4844.get(0);
        mod_4877.put(0, t);
    endrule
    rule rule_6300;
        ChannelMessage t;
        t <- mod_4845.get(1);
        mod_4846.put(0, t);
    endrule
    rule rule_6301;
        ChannelMessage t;
        t <- mod_4845.get(0);
        mod_4870.put(0, t);
    endrule
    rule rule_6302;
        ChannelMessage t;
        t <- mod_4858.get(0);
        mod_4859.put(0, t);
    endrule
    rule rule_6303;
        ChannelMessage t;
        t <- mod_4877.get(0);
        mod_4844.put(1, t);
    endrule
    rule rule_6304;
        ChannelMessage t;
        t <- mod_4862.get(0);
        mod_4850.put(1, t);
    endrule
    rule rule_6305;
        ChannelMessage t;
        t <- mod_4856.get(0);
        mod_4856.put(1, t);
    endrule
    rule rule_6306;
        ChannelMessage t;
        t <- mod_4866.get(1);
        mod_4865.put(1, t);
    endrule
    rule rule_6307;
        ChannelMessage t;
        t <- mod_4841.get(0);
        mod_4842.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_4839.put(0, t);
        end
        if (i == 1) begin
            mod_4855.put(0, t);
        end
        if (i == 2) begin
            mod_4861.put(0, t);
        end
        if (i == 3) begin
            mod_4869.put(0, t);
        end
        if (i == 4) begin
            mod_4875.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 1) begin
            t <- mod_4843.get(0);
        end
        if (i == 0) begin
            t <- mod_4843.get(1);
        end
        if (i == 3) begin
            t <- mod_4843.get(2);
        end
        if (i == 2) begin
            t <- mod_4855.get(0);
        end

        return t;
    endmethod
endmodule

module mkStep(Empty);
    Operation_IFC mod_0_inner <- mkHypernode;
    Operation_IFC mod_0 <- mkDebugOperation(mod_0_inner, "mod_0");
    Operation_IFC mod_41_inner <- mkHypernode;
    Operation_IFC mod_41 <- mkDebugOperation(mod_41_inner, "mod_41");
    Operation_IFC mod_82_inner <- mkHypernode;
    Operation_IFC mod_82 <- mkDebugOperation(mod_82_inner, "mod_82");
    Operation_IFC mod_123_inner <- mkHypernode;
    Operation_IFC mod_123 <- mkDebugOperation(mod_123_inner, "mod_123");
    Operation_IFC mod_164_inner <- mkHypernode;
    Operation_IFC mod_164 <- mkDebugOperation(mod_164_inner, "mod_164");
    Operation_IFC mod_205_inner <- mkHypernode;
    Operation_IFC mod_205 <- mkDebugOperation(mod_205_inner, "mod_205");
    Operation_IFC mod_246_inner <- mkHypernode;
    Operation_IFC mod_246 <- mkDebugOperation(mod_246_inner, "mod_246");
    Operation_IFC mod_287_inner <- mkHypernode;
    Operation_IFC mod_287 <- mkDebugOperation(mod_287_inner, "mod_287");
    Operation_IFC mod_328_inner <- mkHypernode;
    Operation_IFC mod_328 <- mkDebugOperation(mod_328_inner, "mod_328");
    Operation_IFC mod_369_inner <- mkHypernode;
    Operation_IFC mod_369 <- mkDebugOperation(mod_369_inner, "mod_369");
    Operation_IFC mod_410_inner <- mkHypernode;
    Operation_IFC mod_410 <- mkDebugOperation(mod_410_inner, "mod_410");
    Operation_IFC mod_451_inner <- mkHypernode;
    Operation_IFC mod_451 <- mkDebugOperation(mod_451_inner, "mod_451");
    Operation_IFC mod_492_inner <- mkHypernode;
    Operation_IFC mod_492 <- mkDebugOperation(mod_492_inner, "mod_492");
    Operation_IFC mod_533_inner <- mkHypernode;
    Operation_IFC mod_533 <- mkDebugOperation(mod_533_inner, "mod_533");
    Operation_IFC mod_574_inner <- mkHypernode;
    Operation_IFC mod_574 <- mkDebugOperation(mod_574_inner, "mod_574");
    Operation_IFC mod_615_inner <- mkHypernode;
    Operation_IFC mod_615 <- mkDebugOperation(mod_615_inner, "mod_615");
    Operation_IFC mod_656_inner <- mkHypernode;
    Operation_IFC mod_656 <- mkDebugOperation(mod_656_inner, "mod_656");
    Operation_IFC mod_697_inner <- mkHypernode;
    Operation_IFC mod_697 <- mkDebugOperation(mod_697_inner, "mod_697");
    Operation_IFC mod_738_inner <- mkHypernode;
    Operation_IFC mod_738 <- mkDebugOperation(mod_738_inner, "mod_738");
    Operation_IFC mod_779_inner <- mkHypernode;
    Operation_IFC mod_779 <- mkDebugOperation(mod_779_inner, "mod_779");
    Operation_IFC mod_820_inner <- mkHypernode;
    Operation_IFC mod_820 <- mkDebugOperation(mod_820_inner, "mod_820");
    Operation_IFC mod_861_inner <- mkHypernode;
    Operation_IFC mod_861 <- mkDebugOperation(mod_861_inner, "mod_861");
    Operation_IFC mod_902_inner <- mkHypernode;
    Operation_IFC mod_902 <- mkDebugOperation(mod_902_inner, "mod_902");
    Operation_IFC mod_943_inner <- mkHypernode;
    Operation_IFC mod_943 <- mkDebugOperation(mod_943_inner, "mod_943");
    Operation_IFC mod_984_inner <- mkHypernode;
    Operation_IFC mod_984 <- mkDebugOperation(mod_984_inner, "mod_984");
    Operation_IFC mod_1025_inner <- mkHypernode;
    Operation_IFC mod_1025 <- mkDebugOperation(mod_1025_inner, "mod_1025");
    Operation_IFC mod_1066_inner <- mkHypernode;
    Operation_IFC mod_1066 <- mkDebugOperation(mod_1066_inner, "mod_1066");
    Operation_IFC mod_1107_inner <- mkHypernode;
    Operation_IFC mod_1107 <- mkDebugOperation(mod_1107_inner, "mod_1107");
    Operation_IFC mod_1148_inner <- mkHypernode;
    Operation_IFC mod_1148 <- mkDebugOperation(mod_1148_inner, "mod_1148");
    Operation_IFC mod_1189_inner <- mkHypernode;
    Operation_IFC mod_1189 <- mkDebugOperation(mod_1189_inner, "mod_1189");
    Operation_IFC mod_1230_inner <- mkHypernode;
    Operation_IFC mod_1230 <- mkDebugOperation(mod_1230_inner, "mod_1230");
    Operation_IFC mod_1271_inner <- mkHypernode;
    Operation_IFC mod_1271 <- mkDebugOperation(mod_1271_inner, "mod_1271");
    Operation_IFC mod_1312_inner <- mkHypernode;
    Operation_IFC mod_1312 <- mkDebugOperation(mod_1312_inner, "mod_1312");
    Operation_IFC mod_1353_inner <- mkHypernode;
    Operation_IFC mod_1353 <- mkDebugOperation(mod_1353_inner, "mod_1353");
    Operation_IFC mod_1394_inner <- mkHypernode;
    Operation_IFC mod_1394 <- mkDebugOperation(mod_1394_inner, "mod_1394");
    Operation_IFC mod_1435_inner <- mkHypernode;
    Operation_IFC mod_1435 <- mkDebugOperation(mod_1435_inner, "mod_1435");
    Operation_IFC mod_1476_inner <- mkHypernode;
    Operation_IFC mod_1476 <- mkDebugOperation(mod_1476_inner, "mod_1476");
    Operation_IFC mod_1517_inner <- mkHypernode;
    Operation_IFC mod_1517 <- mkDebugOperation(mod_1517_inner, "mod_1517");
    Operation_IFC mod_1558_inner <- mkHypernode;
    Operation_IFC mod_1558 <- mkDebugOperation(mod_1558_inner, "mod_1558");
    Operation_IFC mod_1599_inner <- mkHypernode;
    Operation_IFC mod_1599 <- mkDebugOperation(mod_1599_inner, "mod_1599");
    Operation_IFC mod_1640_inner <- mkHypernode;
    Operation_IFC mod_1640 <- mkDebugOperation(mod_1640_inner, "mod_1640");
    Operation_IFC mod_1681_inner <- mkHypernode;
    Operation_IFC mod_1681 <- mkDebugOperation(mod_1681_inner, "mod_1681");
    Operation_IFC mod_1722_inner <- mkHypernode;
    Operation_IFC mod_1722 <- mkDebugOperation(mod_1722_inner, "mod_1722");
    Operation_IFC mod_1763_inner <- mkHypernode;
    Operation_IFC mod_1763 <- mkDebugOperation(mod_1763_inner, "mod_1763");
    Operation_IFC mod_1804_inner <- mkHypernode;
    Operation_IFC mod_1804 <- mkDebugOperation(mod_1804_inner, "mod_1804");
    Operation_IFC mod_1845_inner <- mkHypernode;
    Operation_IFC mod_1845 <- mkDebugOperation(mod_1845_inner, "mod_1845");
    Operation_IFC mod_1886_inner <- mkHypernode;
    Operation_IFC mod_1886 <- mkDebugOperation(mod_1886_inner, "mod_1886");
    Operation_IFC mod_1927_inner <- mkHypernode;
    Operation_IFC mod_1927 <- mkDebugOperation(mod_1927_inner, "mod_1927");
    Operation_IFC mod_1968_inner <- mkHypernode;
    Operation_IFC mod_1968 <- mkDebugOperation(mod_1968_inner, "mod_1968");
    Operation_IFC mod_2009_inner <- mkHypernode;
    Operation_IFC mod_2009 <- mkDebugOperation(mod_2009_inner, "mod_2009");
    Operation_IFC mod_2050_inner <- mkHypernode;
    Operation_IFC mod_2050 <- mkDebugOperation(mod_2050_inner, "mod_2050");
    Operation_IFC mod_2091_inner <- mkHypernode;
    Operation_IFC mod_2091 <- mkDebugOperation(mod_2091_inner, "mod_2091");
    Operation_IFC mod_2132_inner <- mkHypernode;
    Operation_IFC mod_2132 <- mkDebugOperation(mod_2132_inner, "mod_2132");
    Operation_IFC mod_2173_inner <- mkHypernode;
    Operation_IFC mod_2173 <- mkDebugOperation(mod_2173_inner, "mod_2173");
    Operation_IFC mod_2214_inner <- mkHypernode;
    Operation_IFC mod_2214 <- mkDebugOperation(mod_2214_inner, "mod_2214");
    Operation_IFC mod_2255_inner <- mkHypernode;
    Operation_IFC mod_2255 <- mkDebugOperation(mod_2255_inner, "mod_2255");
    Operation_IFC mod_2296_inner <- mkHypernode;
    Operation_IFC mod_2296 <- mkDebugOperation(mod_2296_inner, "mod_2296");
    Operation_IFC mod_2337_inner <- mkHypernode;
    Operation_IFC mod_2337 <- mkDebugOperation(mod_2337_inner, "mod_2337");
    Operation_IFC mod_2378_inner <- mkHypernode;
    Operation_IFC mod_2378 <- mkDebugOperation(mod_2378_inner, "mod_2378");
    Operation_IFC mod_2419_inner <- mkHypernode;
    Operation_IFC mod_2419 <- mkDebugOperation(mod_2419_inner, "mod_2419");
    Operation_IFC mod_2460_inner <- mkHypernode;
    Operation_IFC mod_2460 <- mkDebugOperation(mod_2460_inner, "mod_2460");
    Operation_IFC mod_2501_inner <- mkHypernode;
    Operation_IFC mod_2501 <- mkDebugOperation(mod_2501_inner, "mod_2501");
    Operation_IFC mod_2542_inner <- mkHypernode;
    Operation_IFC mod_2542 <- mkDebugOperation(mod_2542_inner, "mod_2542");
    Operation_IFC mod_2583_inner <- mkHypernode;
    Operation_IFC mod_2583 <- mkDebugOperation(mod_2583_inner, "mod_2583");
    Operation_IFC mod_2624_inner <- mkHypernode;
    Operation_IFC mod_2624 <- mkDebugOperation(mod_2624_inner, "mod_2624");
    Operation_IFC mod_2665_inner <- mkHypernode;
    Operation_IFC mod_2665 <- mkDebugOperation(mod_2665_inner, "mod_2665");
    Operation_IFC mod_2706_inner <- mkHypernode;
    Operation_IFC mod_2706 <- mkDebugOperation(mod_2706_inner, "mod_2706");
    Operation_IFC mod_2747_inner <- mkHypernode;
    Operation_IFC mod_2747 <- mkDebugOperation(mod_2747_inner, "mod_2747");
    Operation_IFC mod_2788_inner <- mkHypernode;
    Operation_IFC mod_2788 <- mkDebugOperation(mod_2788_inner, "mod_2788");
    Operation_IFC mod_2829_inner <- mkHypernode;
    Operation_IFC mod_2829 <- mkDebugOperation(mod_2829_inner, "mod_2829");
    Operation_IFC mod_2870_inner <- mkHypernode;
    Operation_IFC mod_2870 <- mkDebugOperation(mod_2870_inner, "mod_2870");
    Operation_IFC mod_2911_inner <- mkHypernode;
    Operation_IFC mod_2911 <- mkDebugOperation(mod_2911_inner, "mod_2911");
    Operation_IFC mod_2952_inner <- mkHypernode;
    Operation_IFC mod_2952 <- mkDebugOperation(mod_2952_inner, "mod_2952");
    Operation_IFC mod_2993_inner <- mkHypernode;
    Operation_IFC mod_2993 <- mkDebugOperation(mod_2993_inner, "mod_2993");
    Operation_IFC mod_3034_inner <- mkHypernode;
    Operation_IFC mod_3034 <- mkDebugOperation(mod_3034_inner, "mod_3034");
    Operation_IFC mod_3075_inner <- mkHypernode;
    Operation_IFC mod_3075 <- mkDebugOperation(mod_3075_inner, "mod_3075");
    Operation_IFC mod_3116_inner <- mkHypernode;
    Operation_IFC mod_3116 <- mkDebugOperation(mod_3116_inner, "mod_3116");
    Operation_IFC mod_3157_inner <- mkHypernode;
    Operation_IFC mod_3157 <- mkDebugOperation(mod_3157_inner, "mod_3157");
    Operation_IFC mod_3198_inner <- mkHypernode;
    Operation_IFC mod_3198 <- mkDebugOperation(mod_3198_inner, "mod_3198");
    Operation_IFC mod_3239_inner <- mkHypernode;
    Operation_IFC mod_3239 <- mkDebugOperation(mod_3239_inner, "mod_3239");
    Operation_IFC mod_3280_inner <- mkHypernode;
    Operation_IFC mod_3280 <- mkDebugOperation(mod_3280_inner, "mod_3280");
    Operation_IFC mod_3321_inner <- mkHypernode;
    Operation_IFC mod_3321 <- mkDebugOperation(mod_3321_inner, "mod_3321");
    Operation_IFC mod_3362_inner <- mkHypernode;
    Operation_IFC mod_3362 <- mkDebugOperation(mod_3362_inner, "mod_3362");
    Operation_IFC mod_3403_inner <- mkHypernode;
    Operation_IFC mod_3403 <- mkDebugOperation(mod_3403_inner, "mod_3403");
    Operation_IFC mod_3444_inner <- mkHypernode;
    Operation_IFC mod_3444 <- mkDebugOperation(mod_3444_inner, "mod_3444");
    Operation_IFC mod_3485_inner <- mkHypernode;
    Operation_IFC mod_3485 <- mkDebugOperation(mod_3485_inner, "mod_3485");
    Operation_IFC mod_3526_inner <- mkHypernode;
    Operation_IFC mod_3526 <- mkDebugOperation(mod_3526_inner, "mod_3526");
    Operation_IFC mod_3567_inner <- mkHypernode;
    Operation_IFC mod_3567 <- mkDebugOperation(mod_3567_inner, "mod_3567");
    Operation_IFC mod_3608_inner <- mkHypernode;
    Operation_IFC mod_3608 <- mkDebugOperation(mod_3608_inner, "mod_3608");
    Operation_IFC mod_3649_inner <- mkHypernode;
    Operation_IFC mod_3649 <- mkDebugOperation(mod_3649_inner, "mod_3649");
    Operation_IFC mod_3690_inner <- mkHypernode;
    Operation_IFC mod_3690 <- mkDebugOperation(mod_3690_inner, "mod_3690");
    Operation_IFC mod_3731_inner <- mkHypernode;
    Operation_IFC mod_3731 <- mkDebugOperation(mod_3731_inner, "mod_3731");
    Operation_IFC mod_3772_inner <- mkHypernode;
    Operation_IFC mod_3772 <- mkDebugOperation(mod_3772_inner, "mod_3772");
    Operation_IFC mod_3813_inner <- mkHypernode;
    Operation_IFC mod_3813 <- mkDebugOperation(mod_3813_inner, "mod_3813");
    Operation_IFC mod_3854_inner <- mkHypernode;
    Operation_IFC mod_3854 <- mkDebugOperation(mod_3854_inner, "mod_3854");
    Operation_IFC mod_3895_inner <- mkHypernode;
    Operation_IFC mod_3895 <- mkDebugOperation(mod_3895_inner, "mod_3895");
    Operation_IFC mod_3936_inner <- mkHypernode;
    Operation_IFC mod_3936 <- mkDebugOperation(mod_3936_inner, "mod_3936");
    Operation_IFC mod_3977_inner <- mkHypernode;
    Operation_IFC mod_3977 <- mkDebugOperation(mod_3977_inner, "mod_3977");
    Operation_IFC mod_4018_inner <- mkHypernode;
    Operation_IFC mod_4018 <- mkDebugOperation(mod_4018_inner, "mod_4018");
    Operation_IFC mod_4059_inner <- mkHypernode;
    Operation_IFC mod_4059 <- mkDebugOperation(mod_4059_inner, "mod_4059");
    Operation_IFC mod_4100_inner <- mkHypernode;
    Operation_IFC mod_4100 <- mkDebugOperation(mod_4100_inner, "mod_4100");
    Operation_IFC mod_4141_inner <- mkHypernode;
    Operation_IFC mod_4141 <- mkDebugOperation(mod_4141_inner, "mod_4141");
    Operation_IFC mod_4182_inner <- mkHypernode;
    Operation_IFC mod_4182 <- mkDebugOperation(mod_4182_inner, "mod_4182");
    Operation_IFC mod_4223_inner <- mkHypernode;
    Operation_IFC mod_4223 <- mkDebugOperation(mod_4223_inner, "mod_4223");
    Operation_IFC mod_4264_inner <- mkHypernode;
    Operation_IFC mod_4264 <- mkDebugOperation(mod_4264_inner, "mod_4264");
    Operation_IFC mod_4305_inner <- mkHypernode;
    Operation_IFC mod_4305 <- mkDebugOperation(mod_4305_inner, "mod_4305");
    Operation_IFC mod_4346_inner <- mkHypernode;
    Operation_IFC mod_4346 <- mkDebugOperation(mod_4346_inner, "mod_4346");
    Operation_IFC mod_4387_inner <- mkHypernode;
    Operation_IFC mod_4387 <- mkDebugOperation(mod_4387_inner, "mod_4387");
    Operation_IFC mod_4428_inner <- mkHypernode;
    Operation_IFC mod_4428 <- mkDebugOperation(mod_4428_inner, "mod_4428");
    Operation_IFC mod_4469_inner <- mkHypernode;
    Operation_IFC mod_4469 <- mkDebugOperation(mod_4469_inner, "mod_4469");
    Operation_IFC mod_4510_inner <- mkHypernode;
    Operation_IFC mod_4510 <- mkDebugOperation(mod_4510_inner, "mod_4510");
    Operation_IFC mod_4551_inner <- mkHypernode;
    Operation_IFC mod_4551 <- mkDebugOperation(mod_4551_inner, "mod_4551");
    Operation_IFC mod_4592_inner <- mkHypernode;
    Operation_IFC mod_4592 <- mkDebugOperation(mod_4592_inner, "mod_4592");
    Operation_IFC mod_4633_inner <- mkHypernode;
    Operation_IFC mod_4633 <- mkDebugOperation(mod_4633_inner, "mod_4633");
    Operation_IFC mod_4674_inner <- mkHypernode;
    Operation_IFC mod_4674 <- mkDebugOperation(mod_4674_inner, "mod_4674");
    Operation_IFC mod_4715_inner <- mkHypernode;
    Operation_IFC mod_4715 <- mkDebugOperation(mod_4715_inner, "mod_4715");
    Operation_IFC mod_4756_inner <- mkHypernode;
    Operation_IFC mod_4756 <- mkDebugOperation(mod_4756_inner, "mod_4756");
    Operation_IFC mod_4797_inner <- mkHypernode;
    Operation_IFC mod_4797 <- mkDebugOperation(mod_4797_inner, "mod_4797");
    Operation_IFC mod_4838_inner <- mkHypernode;
    Operation_IFC mod_4838 <- mkDebugOperation(mod_4838_inner, "mod_4838");
    Operation_IFC mod_4879_inner <- mkHypernode;
    Operation_IFC mod_4879 <- mkDebugOperation(mod_4879_inner, "mod_4879");
    Operation_IFC mod_4920_inner <- mkHypernode;
    Operation_IFC mod_4920 <- mkDebugOperation(mod_4920_inner, "mod_4920");
    Operation_IFC mod_4961_inner <- mkHypernode;
    Operation_IFC mod_4961 <- mkDebugOperation(mod_4961_inner, "mod_4961");
    Operation_IFC mod_5002_inner <- mkHypernode;
    Operation_IFC mod_5002 <- mkDebugOperation(mod_5002_inner, "mod_5002");
    Operation_IFC mod_5043_inner <- mkHypernode;
    Operation_IFC mod_5043 <- mkDebugOperation(mod_5043_inner, "mod_5043");
    Operation_IFC mod_5084_inner <- mkHypernode;
    Operation_IFC mod_5084 <- mkDebugOperation(mod_5084_inner, "mod_5084");
    Operation_IFC mod_5125_inner <- mkHypernode;
    Operation_IFC mod_5125 <- mkDebugOperation(mod_5125_inner, "mod_5125");
    Operation_IFC mod_5166_inner <- mkHypernode;
    Operation_IFC mod_5166 <- mkDebugOperation(mod_5166_inner, "mod_5166");
    Operation_IFC mod_5207_inner <- mkHypernode;
    Operation_IFC mod_5207 <- mkDebugOperation(mod_5207_inner, "mod_5207");
    Operation_IFC mod_5248_inner <- mkFlatten(0);
    Operation_IFC mod_5248 <- mkDebugOperation(mod_5248_inner, "mod_5248");
    Operation_IFC mod_5249_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5249 <- mkDebugOperation(mod_5249_inner, "mod_5249");
    Operation_IFC mod_5250_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5250 <- mkDebugOperation(mod_5250_inner, "mod_5250");
    Operation_IFC mod_5251_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5251 <- mkDebugOperation(mod_5251_inner, "mod_5251");
    Operation_IFC mod_5252_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5252 <- mkDebugOperation(mod_5252_inner, "mod_5252");
    Operation_IFC mod_5253_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5253 <- mkDebugOperation(mod_5253_inner, "mod_5253");
    Operation_IFC mod_5254_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5254 <- mkDebugOperation(mod_5254_inner, "mod_5254");
    Operation_IFC mod_5255_inner <- mkPrinter("mod_5255");
    Operation_IFC mod_5255 <- mkDebugOperation(mod_5255_inner, "mod_5255");
    Operation_IFC mod_5256_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5256 <- mkDebugOperation(mod_5256_inner, "mod_5256");
    Operation_IFC mod_5257_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5257 <- mkDebugOperation(mod_5257_inner, "mod_5257");
    Operation_IFC mod_5258_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5258 <- mkDebugOperation(mod_5258_inner, "mod_5258");
    Operation_IFC mod_5259_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5259 <- mkDebugOperation(mod_5259_inner, "mod_5259");
    Operation_IFC mod_5260_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5260 <- mkDebugOperation(mod_5260_inner, "mod_5260");
    Operation_IFC mod_5261_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5261 <- mkDebugOperation(mod_5261_inner, "mod_5261");
    Operation_IFC mod_5262_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5262 <- mkDebugOperation(mod_5262_inner, "mod_5262");
    Operation_IFC mod_5263_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5263 <- mkDebugOperation(mod_5263_inner, "mod_5263");
    Operation_IFC mod_5264_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5264 <- mkDebugOperation(mod_5264_inner, "mod_5264");
    Operation_IFC mod_5265_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5265 <- mkDebugOperation(mod_5265_inner, "mod_5265");
    Operation_IFC mod_5266_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5266 <- mkDebugOperation(mod_5266_inner, "mod_5266");
    Operation_IFC mod_5267_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5267 <- mkDebugOperation(mod_5267_inner, "mod_5267");
    Operation_IFC mod_5268_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5268 <- mkDebugOperation(mod_5268_inner, "mod_5268");
    Operation_IFC mod_5269_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5269 <- mkDebugOperation(mod_5269_inner, "mod_5269");
    Operation_IFC mod_5270_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5270 <- mkDebugOperation(mod_5270_inner, "mod_5270");
    Operation_IFC mod_5271_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5271 <- mkDebugOperation(mod_5271_inner, "mod_5271");
    Operation_IFC mod_5272_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5272 <- mkDebugOperation(mod_5272_inner, "mod_5272");
    Operation_IFC mod_5273_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5273 <- mkDebugOperation(mod_5273_inner, "mod_5273");
    Operation_IFC mod_5274_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5274 <- mkDebugOperation(mod_5274_inner, "mod_5274");
    Operation_IFC mod_5275_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5275 <- mkDebugOperation(mod_5275_inner, "mod_5275");
    Operation_IFC mod_5276_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5276 <- mkDebugOperation(mod_5276_inner, "mod_5276");
    Operation_IFC mod_5277_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5277 <- mkDebugOperation(mod_5277_inner, "mod_5277");
    Operation_IFC mod_5278_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5278 <- mkDebugOperation(mod_5278_inner, "mod_5278");
    Operation_IFC mod_5279_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5279 <- mkDebugOperation(mod_5279_inner, "mod_5279");
    Operation_IFC mod_5280_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5280 <- mkDebugOperation(mod_5280_inner, "mod_5280");
    Operation_IFC mod_5281_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5281 <- mkDebugOperation(mod_5281_inner, "mod_5281");
    Operation_IFC mod_5282_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5282 <- mkDebugOperation(mod_5282_inner, "mod_5282");
    Operation_IFC mod_5283_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5283 <- mkDebugOperation(mod_5283_inner, "mod_5283");
    Operation_IFC mod_5284_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5284 <- mkDebugOperation(mod_5284_inner, "mod_5284");
    Operation_IFC mod_5285_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5285 <- mkDebugOperation(mod_5285_inner, "mod_5285");
    Operation_IFC mod_5286_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5286 <- mkDebugOperation(mod_5286_inner, "mod_5286");
    Operation_IFC mod_5287_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5287 <- mkDebugOperation(mod_5287_inner, "mod_5287");
    Operation_IFC mod_5288_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5288 <- mkDebugOperation(mod_5288_inner, "mod_5288");
    Operation_IFC mod_5289_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5289 <- mkDebugOperation(mod_5289_inner, "mod_5289");
    Operation_IFC mod_5290_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5290 <- mkDebugOperation(mod_5290_inner, "mod_5290");
    Operation_IFC mod_5291_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5291 <- mkDebugOperation(mod_5291_inner, "mod_5291");
    Operation_IFC mod_5292_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5292 <- mkDebugOperation(mod_5292_inner, "mod_5292");
    Operation_IFC mod_5293_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5293 <- mkDebugOperation(mod_5293_inner, "mod_5293");
    Operation_IFC mod_5294_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5294 <- mkDebugOperation(mod_5294_inner, "mod_5294");
    Operation_IFC mod_5295_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5295 <- mkDebugOperation(mod_5295_inner, "mod_5295");
    Operation_IFC mod_5296_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5296 <- mkDebugOperation(mod_5296_inner, "mod_5296");
    Operation_IFC mod_5297_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5297 <- mkDebugOperation(mod_5297_inner, "mod_5297");
    Operation_IFC mod_5298_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5298 <- mkDebugOperation(mod_5298_inner, "mod_5298");
    Operation_IFC mod_5299_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5299 <- mkDebugOperation(mod_5299_inner, "mod_5299");
    Operation_IFC mod_5300_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5300 <- mkDebugOperation(mod_5300_inner, "mod_5300");
    Operation_IFC mod_5301_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5301 <- mkDebugOperation(mod_5301_inner, "mod_5301");
    Operation_IFC mod_5302_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5302 <- mkDebugOperation(mod_5302_inner, "mod_5302");
    Operation_IFC mod_5303_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5303 <- mkDebugOperation(mod_5303_inner, "mod_5303");
    Operation_IFC mod_5304_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5304 <- mkDebugOperation(mod_5304_inner, "mod_5304");
    Operation_IFC mod_5305_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5305 <- mkDebugOperation(mod_5305_inner, "mod_5305");
    Operation_IFC mod_5306_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5306 <- mkDebugOperation(mod_5306_inner, "mod_5306");
    Operation_IFC mod_5307_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5307 <- mkDebugOperation(mod_5307_inner, "mod_5307");
    Operation_IFC mod_5308_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5308 <- mkDebugOperation(mod_5308_inner, "mod_5308");
    Partition_IFC#(128) mod_5309_inner <- mkPartition(0, 128);
    Operation_IFC mod_5309 <- mkDebugOperation(mod_5309_inner.op, "mod_5309");
    Operation_IFC mod_5310_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5310 <- mkDebugOperation(mod_5310_inner, "mod_5310");
    Operation_IFC mod_5311_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5311 <- mkDebugOperation(mod_5311_inner, "mod_5311");
    Operation_IFC mod_5312_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5312 <- mkDebugOperation(mod_5312_inner, "mod_5312");
    Reassemble_IFC#(128) mod_5313_inner <- mkReassemble(128);
    Operation_IFC mod_5313 <- mkDebugOperation(mod_5313_inner.op, "mod_5313");
    Operation_IFC mod_5314_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5314 <- mkDebugOperation(mod_5314_inner, "mod_5314");
    Operation_IFC mod_5315_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5315 <- mkDebugOperation(mod_5315_inner, "mod_5315");
    Operation_IFC mod_5316_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5316 <- mkDebugOperation(mod_5316_inner, "mod_5316");
    Operation_IFC mod_5317_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5317 <- mkDebugOperation(mod_5317_inner, "mod_5317");
    Operation_IFC mod_5318_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5318 <- mkDebugOperation(mod_5318_inner, "mod_5318");
    Operation_IFC mod_5319_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5319 <- mkDebugOperation(mod_5319_inner, "mod_5319");
    Operation_IFC mod_5320_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5320 <- mkDebugOperation(mod_5320_inner, "mod_5320");
    Operation_IFC mod_5321_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5321 <- mkDebugOperation(mod_5321_inner, "mod_5321");
    Operation_IFC mod_5322_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5322 <- mkDebugOperation(mod_5322_inner, "mod_5322");
    Operation_IFC mod_5323_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5323 <- mkDebugOperation(mod_5323_inner, "mod_5323");
    Operation_IFC mod_5324_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5324 <- mkDebugOperation(mod_5324_inner, "mod_5324");
    Operation_IFC mod_5325_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5325 <- mkDebugOperation(mod_5325_inner, "mod_5325");
    PMU_IFC mod_5326_bufferize <- mkPMU(2);
    Operation_IFC mod_5326_inner = mod_5326_bufferize.operation;
    Operation_IFC mod_5326 <- mkDebugOperation(mod_5326_inner, "mod_5326");
    Operation_IFC mod_5327_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5327 <- mkDebugOperation(mod_5327_inner, "mod_5327");
    Operation_IFC mod_5328_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5328 <- mkDebugOperation(mod_5328_inner, "mod_5328");
    Operation_IFC mod_5329_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5329 <- mkDebugOperation(mod_5329_inner, "mod_5329");
    Operation_IFC mod_5330_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5330 <- mkDebugOperation(mod_5330_inner, "mod_5330");
    Operation_IFC mod_5331_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5331 <- mkDebugOperation(mod_5331_inner, "mod_5331");
    Operation_IFC mod_5332_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5332 <- mkDebugOperation(mod_5332_inner, "mod_5332");
    Operation_IFC mod_5333_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5333 <- mkDebugOperation(mod_5333_inner, "mod_5333");
    Operation_IFC mod_5334_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5334 <- mkDebugOperation(mod_5334_inner, "mod_5334");
    Operation_IFC mod_5335_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5335 <- mkDebugOperation(mod_5335_inner, "mod_5335");
    Operation_IFC mod_5336_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5336 <- mkDebugOperation(mod_5336_inner, "mod_5336");
    Operation_IFC mod_5337_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5337 <- mkDebugOperation(mod_5337_inner, "mod_5337");
    Operation_IFC mod_5338_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5338 <- mkDebugOperation(mod_5338_inner, "mod_5338");
    Operation_IFC mod_5339_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5339 <- mkDebugOperation(mod_5339_inner, "mod_5339");
    Operation_IFC mod_5340_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5340 <- mkDebugOperation(mod_5340_inner, "mod_5340");
    Operation_IFC mod_5341_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5341 <- mkDebugOperation(mod_5341_inner, "mod_5341");
    Operation_IFC mod_5342_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5342 <- mkDebugOperation(mod_5342_inner, "mod_5342");
    Operation_IFC mod_5343_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5343 <- mkDebugOperation(mod_5343_inner, "mod_5343");
    Operation_IFC mod_5344_inner <- mkRandomOffChipLoad(Cons(64, Cons(1, Cons(1, Cons(1, Cons(1, Cons(1, Nil)))))));
    Operation_IFC mod_5344 <- mkDebugOperation(mod_5344_inner, "mod_5344");
    Operation_IFC mod_5345_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5345 <- mkDebugOperation(mod_5345_inner, "mod_5345");
    Operation_IFC mod_5346_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5346 <- mkDebugOperation(mod_5346_inner, "mod_5346");
    Operation_IFC mod_5347_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5347 <- mkDebugOperation(mod_5347_inner, "mod_5347");
    Operation_IFC mod_5348_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5348 <- mkDebugOperation(mod_5348_inner, "mod_5348");
    Operation_IFC mod_5349_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5349 <- mkDebugOperation(mod_5349_inner, "mod_5349");
    Operation_IFC mod_5350_inner <- mkRandomSelectGen(128);
    Operation_IFC mod_5350 <- mkDebugOperation(mod_5350_inner, "mod_5350");
    Operation_IFC mod_5351_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5351 <- mkDebugOperation(mod_5351_inner, "mod_5351");
    Operation_IFC mod_5352_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5352 <- mkDebugOperation(mod_5352_inner, "mod_5352");
    Operation_IFC mod_5353_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5353 <- mkDebugOperation(mod_5353_inner, "mod_5353");
    Operation_IFC mod_5354_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5354 <- mkDebugOperation(mod_5354_inner, "mod_5354");
    Operation_IFC mod_5355_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5355 <- mkDebugOperation(mod_5355_inner, "mod_5355");
    Operation_IFC mod_5356_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5356 <- mkDebugOperation(mod_5356_inner, "mod_5356");
    Operation_IFC mod_5357_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5357 <- mkDebugOperation(mod_5357_inner, "mod_5357");
    Operation_IFC mod_5358_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5358 <- mkDebugOperation(mod_5358_inner, "mod_5358");
    Operation_IFC mod_5359_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5359 <- mkDebugOperation(mod_5359_inner, "mod_5359");
    Operation_IFC mod_5360_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5360 <- mkDebugOperation(mod_5360_inner, "mod_5360");
    Operation_IFC mod_5361_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5361 <- mkDebugOperation(mod_5361_inner, "mod_5361");
    Operation_IFC mod_5362_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5362 <- mkDebugOperation(mod_5362_inner, "mod_5362");
    Operation_IFC mod_5363_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5363 <- mkDebugOperation(mod_5363_inner, "mod_5363");
    Operation_IFC mod_5364_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5364 <- mkDebugOperation(mod_5364_inner, "mod_5364");
    Operation_IFC mod_5365_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5365 <- mkDebugOperation(mod_5365_inner, "mod_5365");
    Operation_IFC mod_5366_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5366 <- mkDebugOperation(mod_5366_inner, "mod_5366");
    Operation_IFC mod_5367_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5367 <- mkDebugOperation(mod_5367_inner, "mod_5367");
    Operation_IFC mod_5368_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5368 <- mkDebugOperation(mod_5368_inner, "mod_5368");
    Operation_IFC mod_5369_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5369 <- mkDebugOperation(mod_5369_inner, "mod_5369");
    Operation_IFC mod_5370_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5370 <- mkDebugOperation(mod_5370_inner, "mod_5370");
    Operation_IFC mod_5371_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5371 <- mkDebugOperation(mod_5371_inner, "mod_5371");
    Operation_IFC mod_5372_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_5372 <- mkDebugOperation(mod_5372_inner, "mod_5372");
    Operation_IFC mod_5373_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5373 <- mkDebugOperation(mod_5373_inner, "mod_5373");
    Operation_IFC mod_5374_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5374 <- mkDebugOperation(mod_5374_inner, "mod_5374");
    Operation_IFC mod_5375_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5375 <- mkDebugOperation(mod_5375_inner, "mod_5375");
    Operation_IFC mod_5376_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5376 <- mkDebugOperation(mod_5376_inner, "mod_5376");
    Operation_IFC mod_5377_inner <- mkRepeatStatic(1);
    Operation_IFC mod_5377 <- mkDebugOperation(mod_5377_inner, "mod_5377");
    Operation_IFC mod_5378_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5378 <- mkDebugOperation(mod_5378_inner, "mod_5378");
    Operation_IFC mod_5379_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5379 <- mkDebugOperation(mod_5379_inner, "mod_5379");
    Operation_IFC mod_5380_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5380 <- mkDebugOperation(mod_5380_inner, "mod_5380");
    Operation_IFC mod_5381_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5381 <- mkDebugOperation(mod_5381_inner, "mod_5381");
    Operation_IFC mod_5382_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5382 <- mkDebugOperation(mod_5382_inner, "mod_5382");
    Operation_IFC mod_5383_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5383 <- mkDebugOperation(mod_5383_inner, "mod_5383");
    Operation_IFC mod_5384_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5384 <- mkDebugOperation(mod_5384_inner, "mod_5384");
    Operation_IFC mod_5385_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5385 <- mkDebugOperation(mod_5385_inner, "mod_5385");
    Operation_IFC mod_5386_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5386 <- mkDebugOperation(mod_5386_inner, "mod_5386");
    Operation_IFC mod_5387_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5387 <- mkDebugOperation(mod_5387_inner, "mod_5387");
    Operation_IFC mod_5388_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5388 <- mkDebugOperation(mod_5388_inner, "mod_5388");
    Operation_IFC mod_5389_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5389 <- mkDebugOperation(mod_5389_inner, "mod_5389");
    Operation_IFC mod_5390_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5390 <- mkDebugOperation(mod_5390_inner, "mod_5390");
    Operation_IFC mod_5391_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5391 <- mkDebugOperation(mod_5391_inner, "mod_5391");
    Operation_IFC mod_5392_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5392 <- mkDebugOperation(mod_5392_inner, "mod_5392");
    Operation_IFC mod_5393_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5393 <- mkDebugOperation(mod_5393_inner, "mod_5393");
    Operation_IFC mod_5394_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5394 <- mkDebugOperation(mod_5394_inner, "mod_5394");
    Operation_IFC mod_5395_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5395 <- mkDebugOperation(mod_5395_inner, "mod_5395");
    Operation_IFC mod_5396_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5396 <- mkDebugOperation(mod_5396_inner, "mod_5396");
    Operation_IFC mod_5397_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5397 <- mkDebugOperation(mod_5397_inner, "mod_5397");
    Operation_IFC mod_5398_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5398 <- mkDebugOperation(mod_5398_inner, "mod_5398");
    Operation_IFC mod_5399_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5399 <- mkDebugOperation(mod_5399_inner, "mod_5399");
    Operation_IFC mod_5400_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5400 <- mkDebugOperation(mod_5400_inner, "mod_5400");
    Operation_IFC mod_5401_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5401 <- mkDebugOperation(mod_5401_inner, "mod_5401");
    Operation_IFC mod_5402_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5402 <- mkDebugOperation(mod_5402_inner, "mod_5402");
    Operation_IFC mod_5403_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5403 <- mkDebugOperation(mod_5403_inner, "mod_5403");
    Operation_IFC mod_5404_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5404 <- mkDebugOperation(mod_5404_inner, "mod_5404");
    Operation_IFC mod_5405_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5405 <- mkDebugOperation(mod_5405_inner, "mod_5405");
    Operation_IFC mod_5406_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5406 <- mkDebugOperation(mod_5406_inner, "mod_5406");
    Operation_IFC mod_5407_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5407 <- mkDebugOperation(mod_5407_inner, "mod_5407");
    Operation_IFC mod_5408_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5408 <- mkDebugOperation(mod_5408_inner, "mod_5408");
    Operation_IFC mod_5409_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5409 <- mkDebugOperation(mod_5409_inner, "mod_5409");
    Operation_IFC mod_5410_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5410 <- mkDebugOperation(mod_5410_inner, "mod_5410");
    Operation_IFC mod_5411_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5411 <- mkDebugOperation(mod_5411_inner, "mod_5411");
    Operation_IFC mod_5412_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5412 <- mkDebugOperation(mod_5412_inner, "mod_5412");
    Operation_IFC mod_5413_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5413 <- mkDebugOperation(mod_5413_inner, "mod_5413");
    Operation_IFC mod_5414_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5414 <- mkDebugOperation(mod_5414_inner, "mod_5414");
    Operation_IFC mod_5415_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5415 <- mkDebugOperation(mod_5415_inner, "mod_5415");
    Operation_IFC mod_5416_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5416 <- mkDebugOperation(mod_5416_inner, "mod_5416");
    Operation_IFC mod_5417_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5417 <- mkDebugOperation(mod_5417_inner, "mod_5417");
    Operation_IFC mod_5418_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5418 <- mkDebugOperation(mod_5418_inner, "mod_5418");
    Operation_IFC mod_5419_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5419 <- mkDebugOperation(mod_5419_inner, "mod_5419");
    Operation_IFC mod_5420_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5420 <- mkDebugOperation(mod_5420_inner, "mod_5420");
    Operation_IFC mod_5421_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5421 <- mkDebugOperation(mod_5421_inner, "mod_5421");
    Operation_IFC mod_5422_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5422 <- mkDebugOperation(mod_5422_inner, "mod_5422");
    Operation_IFC mod_5423_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5423 <- mkDebugOperation(mod_5423_inner, "mod_5423");
    Operation_IFC mod_5424_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5424 <- mkDebugOperation(mod_5424_inner, "mod_5424");
    Operation_IFC mod_5425_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5425 <- mkDebugOperation(mod_5425_inner, "mod_5425");
    Operation_IFC mod_5426_inner <- mkRandomSelectGen(128);
    Operation_IFC mod_5426 <- mkDebugOperation(mod_5426_inner, "mod_5426");
    Operation_IFC mod_5427_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5427 <- mkDebugOperation(mod_5427_inner, "mod_5427");
    Operation_IFC mod_5428_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5428 <- mkDebugOperation(mod_5428_inner, "mod_5428");
    Operation_IFC mod_5429_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5429 <- mkDebugOperation(mod_5429_inner, "mod_5429");
    Operation_IFC mod_5430_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5430 <- mkDebugOperation(mod_5430_inner, "mod_5430");
    Operation_IFC mod_5431_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5431 <- mkDebugOperation(mod_5431_inner, "mod_5431");
    Operation_IFC mod_5432_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5432 <- mkDebugOperation(mod_5432_inner, "mod_5432");
    Operation_IFC mod_5433_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5433 <- mkDebugOperation(mod_5433_inner, "mod_5433");
    Operation_IFC mod_5434_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5434 <- mkDebugOperation(mod_5434_inner, "mod_5434");
    Operation_IFC mod_5435_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5435 <- mkDebugOperation(mod_5435_inner, "mod_5435");
    Operation_IFC mod_5436_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5436 <- mkDebugOperation(mod_5436_inner, "mod_5436");
    Operation_IFC mod_5437_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5437 <- mkDebugOperation(mod_5437_inner, "mod_5437");
    Operation_IFC mod_5438_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5438 <- mkDebugOperation(mod_5438_inner, "mod_5438");
    Operation_IFC mod_5439_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5439 <- mkDebugOperation(mod_5439_inner, "mod_5439");
    Operation_IFC mod_5440_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5440 <- mkDebugOperation(mod_5440_inner, "mod_5440");
    Operation_IFC mod_5441_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5441 <- mkDebugOperation(mod_5441_inner, "mod_5441");
    Operation_IFC mod_5442_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5442 <- mkDebugOperation(mod_5442_inner, "mod_5442");
    Operation_IFC mod_5443_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5443 <- mkDebugOperation(mod_5443_inner, "mod_5443");
    Operation_IFC mod_5444_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5444 <- mkDebugOperation(mod_5444_inner, "mod_5444");
    Operation_IFC mod_5445_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5445 <- mkDebugOperation(mod_5445_inner, "mod_5445");
    Operation_IFC mod_5446_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5446 <- mkDebugOperation(mod_5446_inner, "mod_5446");
    Operation_IFC mod_5447_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5447 <- mkDebugOperation(mod_5447_inner, "mod_5447");
    Operation_IFC mod_5448_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5448 <- mkDebugOperation(mod_5448_inner, "mod_5448");
    Operation_IFC mod_5449_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5449 <- mkDebugOperation(mod_5449_inner, "mod_5449");
    Operation_IFC mod_5450_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5450 <- mkDebugOperation(mod_5450_inner, "mod_5450");
    Operation_IFC mod_5451_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5451 <- mkDebugOperation(mod_5451_inner, "mod_5451");
    Operation_IFC mod_5452_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5452 <- mkDebugOperation(mod_5452_inner, "mod_5452");
    Operation_IFC mod_5453_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5453 <- mkDebugOperation(mod_5453_inner, "mod_5453");
    Operation_IFC mod_5454_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5454 <- mkDebugOperation(mod_5454_inner, "mod_5454");
    Operation_IFC mod_5455_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5455 <- mkDebugOperation(mod_5455_inner, "mod_5455");
    Operation_IFC mod_5456_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5456 <- mkDebugOperation(mod_5456_inner, "mod_5456");
    Operation_IFC mod_5457_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5457 <- mkDebugOperation(mod_5457_inner, "mod_5457");
    Operation_IFC mod_5458_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5458 <- mkDebugOperation(mod_5458_inner, "mod_5458");
    Operation_IFC mod_5459_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5459 <- mkDebugOperation(mod_5459_inner, "mod_5459");
    Operation_IFC mod_5460_inner <- mkRandomOffChipLoad(Cons(64, Cons(8, Cons(1, Cons(1, Cons(1, Cons(1, Nil)))))));
    Operation_IFC mod_5460 <- mkDebugOperation(mod_5460_inner, "mod_5460");
    Operation_IFC mod_5461_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5461 <- mkDebugOperation(mod_5461_inner, "mod_5461");
    Operation_IFC mod_5462_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5462 <- mkDebugOperation(mod_5462_inner, "mod_5462");
    Operation_IFC mod_5463_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5463 <- mkDebugOperation(mod_5463_inner, "mod_5463");
    Operation_IFC mod_5464_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5464 <- mkDebugOperation(mod_5464_inner, "mod_5464");
    Operation_IFC mod_5465_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5465 <- mkDebugOperation(mod_5465_inner, "mod_5465");
    Operation_IFC mod_5466_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5466 <- mkDebugOperation(mod_5466_inner, "mod_5466");
    Operation_IFC mod_5467_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5467 <- mkDebugOperation(mod_5467_inner, "mod_5467");
    Operation_IFC mod_5468_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5468 <- mkDebugOperation(mod_5468_inner, "mod_5468");
    Operation_IFC mod_5469_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5469 <- mkDebugOperation(mod_5469_inner, "mod_5469");
    Operation_IFC mod_5470_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5470 <- mkDebugOperation(mod_5470_inner, "mod_5470");
    Operation_IFC mod_5471_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5471 <- mkDebugOperation(mod_5471_inner, "mod_5471");
    Operation_IFC mod_5472_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5472 <- mkDebugOperation(mod_5472_inner, "mod_5472");
    Operation_IFC mod_5473_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5473 <- mkDebugOperation(mod_5473_inner, "mod_5473");
    Operation_IFC mod_5474_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5474 <- mkDebugOperation(mod_5474_inner, "mod_5474");
    Operation_IFC mod_5475_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5475 <- mkDebugOperation(mod_5475_inner, "mod_5475");
    Operation_IFC mod_5476_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5476 <- mkDebugOperation(mod_5476_inner, "mod_5476");
    Operation_IFC mod_5477_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5477 <- mkDebugOperation(mod_5477_inner, "mod_5477");
    Operation_IFC mod_5478_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5478 <- mkDebugOperation(mod_5478_inner, "mod_5478");
    Operation_IFC mod_5479_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5479 <- mkDebugOperation(mod_5479_inner, "mod_5479");
    Operation_IFC mod_5480_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5480 <- mkDebugOperation(mod_5480_inner, "mod_5480");
    Operation_IFC mod_5481_inner <- mkRandomSelectGen(128);
    Operation_IFC mod_5481 <- mkDebugOperation(mod_5481_inner, "mod_5481");
    Operation_IFC mod_5482_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5482 <- mkDebugOperation(mod_5482_inner, "mod_5482");
    Operation_IFC mod_5483_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5483 <- mkDebugOperation(mod_5483_inner, "mod_5483");
    Operation_IFC mod_5484_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5484 <- mkDebugOperation(mod_5484_inner, "mod_5484");
    Operation_IFC mod_5485_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5485 <- mkDebugOperation(mod_5485_inner, "mod_5485");
    Operation_IFC mod_5486_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5486 <- mkDebugOperation(mod_5486_inner, "mod_5486");
    Operation_IFC mod_5487_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5487 <- mkDebugOperation(mod_5487_inner, "mod_5487");
    Operation_IFC mod_5488_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5488 <- mkDebugOperation(mod_5488_inner, "mod_5488");
    Operation_IFC mod_5489_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5489 <- mkDebugOperation(mod_5489_inner, "mod_5489");
    Operation_IFC mod_5490_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5490 <- mkDebugOperation(mod_5490_inner, "mod_5490");
    Operation_IFC mod_5491_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5491 <- mkDebugOperation(mod_5491_inner, "mod_5491");
    Operation_IFC mod_5492_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5492 <- mkDebugOperation(mod_5492_inner, "mod_5492");
    Operation_IFC mod_5493_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5493 <- mkDebugOperation(mod_5493_inner, "mod_5493");
    Operation_IFC mod_5494_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5494 <- mkDebugOperation(mod_5494_inner, "mod_5494");
    Operation_IFC mod_5495_inner <- mkReshape(2, 1);
    Operation_IFC mod_5495 <- mkDebugOperation(mod_5495_inner, "mod_5495");
    Operation_IFC mod_5496_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5496 <- mkDebugOperation(mod_5496_inner, "mod_5496");
    Operation_IFC mod_5497_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5497 <- mkDebugOperation(mod_5497_inner, "mod_5497");
    Operation_IFC mod_5498_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5498 <- mkDebugOperation(mod_5498_inner, "mod_5498");
    Operation_IFC mod_5499_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5499 <- mkDebugOperation(mod_5499_inner, "mod_5499");
    Operation_IFC mod_5500_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5500 <- mkDebugOperation(mod_5500_inner, "mod_5500");
    Operation_IFC mod_5501_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5501 <- mkDebugOperation(mod_5501_inner, "mod_5501");
    Operation_IFC mod_5502_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5502 <- mkDebugOperation(mod_5502_inner, "mod_5502");
    Operation_IFC mod_5503_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5503 <- mkDebugOperation(mod_5503_inner, "mod_5503");
    Operation_IFC mod_5504_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5504 <- mkDebugOperation(mod_5504_inner, "mod_5504");
    Operation_IFC mod_5505_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5505 <- mkDebugOperation(mod_5505_inner, "mod_5505");
    Operation_IFC mod_5506_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5506 <- mkDebugOperation(mod_5506_inner, "mod_5506");
    Operation_IFC mod_5507_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5507 <- mkDebugOperation(mod_5507_inner, "mod_5507");
    Operation_IFC mod_5508_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5508 <- mkDebugOperation(mod_5508_inner, "mod_5508");
    Operation_IFC mod_5509_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5509 <- mkDebugOperation(mod_5509_inner, "mod_5509");
    Operation_IFC mod_5510_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5510 <- mkDebugOperation(mod_5510_inner, "mod_5510");
    Operation_IFC mod_5511_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5511 <- mkDebugOperation(mod_5511_inner, "mod_5511");
    Operation_IFC mod_5512_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5512 <- mkDebugOperation(mod_5512_inner, "mod_5512");
    Operation_IFC mod_5513_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5513 <- mkDebugOperation(mod_5513_inner, "mod_5513");
    Operation_IFC mod_5514_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5514 <- mkDebugOperation(mod_5514_inner, "mod_5514");
    Operation_IFC mod_5515_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5515 <- mkDebugOperation(mod_5515_inner, "mod_5515");
    Operation_IFC mod_5516_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5516 <- mkDebugOperation(mod_5516_inner, "mod_5516");
    Operation_IFC mod_5517_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5517 <- mkDebugOperation(mod_5517_inner, "mod_5517");
    Operation_IFC mod_5518_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5518 <- mkDebugOperation(mod_5518_inner, "mod_5518");
    Operation_IFC mod_5519_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5519 <- mkDebugOperation(mod_5519_inner, "mod_5519");
    Operation_IFC mod_5520_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5520 <- mkDebugOperation(mod_5520_inner, "mod_5520");
    Operation_IFC mod_5521_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5521 <- mkDebugOperation(mod_5521_inner, "mod_5521");
    Operation_IFC mod_5522_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5522 <- mkDebugOperation(mod_5522_inner, "mod_5522");
    Operation_IFC mod_5523_inner <- mkRepeatStatic(1);
    Operation_IFC mod_5523 <- mkDebugOperation(mod_5523_inner, "mod_5523");
    Operation_IFC mod_5524_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5524 <- mkDebugOperation(mod_5524_inner, "mod_5524");
    Operation_IFC mod_5525_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5525 <- mkDebugOperation(mod_5525_inner, "mod_5525");
    Operation_IFC mod_5526_inner <- mkRepeatStatic(1);
    Operation_IFC mod_5526 <- mkDebugOperation(mod_5526_inner, "mod_5526");
    Operation_IFC mod_5527_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5527 <- mkDebugOperation(mod_5527_inner, "mod_5527");
    Operation_IFC mod_5528_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5528 <- mkDebugOperation(mod_5528_inner, "mod_5528");
    Operation_IFC mod_5529_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5529 <- mkDebugOperation(mod_5529_inner, "mod_5529");
    Operation_IFC mod_5530_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5530 <- mkDebugOperation(mod_5530_inner, "mod_5530");
    Operation_IFC mod_5531_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5531 <- mkDebugOperation(mod_5531_inner, "mod_5531");
    Operation_IFC mod_5532_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5532 <- mkDebugOperation(mod_5532_inner, "mod_5532");
    Operation_IFC mod_5533_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5533 <- mkDebugOperation(mod_5533_inner, "mod_5533");
    Operation_IFC mod_5534_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5534 <- mkDebugOperation(mod_5534_inner, "mod_5534");
    Operation_IFC mod_5535_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5535 <- mkDebugOperation(mod_5535_inner, "mod_5535");
    Operation_IFC mod_5536_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5536 <- mkDebugOperation(mod_5536_inner, "mod_5536");
    Operation_IFC mod_5537_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5537 <- mkDebugOperation(mod_5537_inner, "mod_5537");
    Operation_IFC mod_5538_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5538 <- mkDebugOperation(mod_5538_inner, "mod_5538");
    Operation_IFC mod_5539_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5539 <- mkDebugOperation(mod_5539_inner, "mod_5539");
    Operation_IFC mod_5540_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5540 <- mkDebugOperation(mod_5540_inner, "mod_5540");
    Operation_IFC mod_5541_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5541 <- mkDebugOperation(mod_5541_inner, "mod_5541");
    Operation_IFC mod_5542_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5542 <- mkDebugOperation(mod_5542_inner, "mod_5542");
    Operation_IFC mod_5543_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5543 <- mkDebugOperation(mod_5543_inner, "mod_5543");
    Operation_IFC mod_5544_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5544 <- mkDebugOperation(mod_5544_inner, "mod_5544");
    Operation_IFC mod_5545_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5545 <- mkDebugOperation(mod_5545_inner, "mod_5545");
    Operation_IFC mod_5546_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5546 <- mkDebugOperation(mod_5546_inner, "mod_5546");
    Operation_IFC mod_5547_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5547 <- mkDebugOperation(mod_5547_inner, "mod_5547");
    Operation_IFC mod_5548_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5548 <- mkDebugOperation(mod_5548_inner, "mod_5548");
    Operation_IFC mod_5549_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5549 <- mkDebugOperation(mod_5549_inner, "mod_5549");
    Operation_IFC mod_5550_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5550 <- mkDebugOperation(mod_5550_inner, "mod_5550");
    Operation_IFC mod_5551_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5551 <- mkDebugOperation(mod_5551_inner, "mod_5551");
    Operation_IFC mod_5552_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5552 <- mkDebugOperation(mod_5552_inner, "mod_5552");
    Operation_IFC mod_5553_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5553 <- mkDebugOperation(mod_5553_inner, "mod_5553");
    Operation_IFC mod_5554_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5554 <- mkDebugOperation(mod_5554_inner, "mod_5554");
    Operation_IFC mod_5555_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5555 <- mkDebugOperation(mod_5555_inner, "mod_5555");
    Operation_IFC mod_5556_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5556 <- mkDebugOperation(mod_5556_inner, "mod_5556");
    Operation_IFC mod_5557_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5557 <- mkDebugOperation(mod_5557_inner, "mod_5557");
    Operation_IFC mod_5558_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5558 <- mkDebugOperation(mod_5558_inner, "mod_5558");
    Operation_IFC mod_5559_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5559 <- mkDebugOperation(mod_5559_inner, "mod_5559");
    Operation_IFC mod_5560_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5560 <- mkDebugOperation(mod_5560_inner, "mod_5560");
    Operation_IFC mod_5561_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5561 <- mkDebugOperation(mod_5561_inner, "mod_5561");
    Operation_IFC mod_5562_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5562 <- mkDebugOperation(mod_5562_inner, "mod_5562");
    Operation_IFC mod_5563_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5563 <- mkDebugOperation(mod_5563_inner, "mod_5563");
    Operation_IFC mod_5564_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5564 <- mkDebugOperation(mod_5564_inner, "mod_5564");
    Operation_IFC mod_5565_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5565 <- mkDebugOperation(mod_5565_inner, "mod_5565");
    Operation_IFC mod_5566_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5566 <- mkDebugOperation(mod_5566_inner, "mod_5566");
    Operation_IFC mod_5567_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5567 <- mkDebugOperation(mod_5567_inner, "mod_5567");
    Operation_IFC mod_5568_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5568 <- mkDebugOperation(mod_5568_inner, "mod_5568");
    Operation_IFC mod_5569_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5569 <- mkDebugOperation(mod_5569_inner, "mod_5569");
    Operation_IFC mod_5570_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5570 <- mkDebugOperation(mod_5570_inner, "mod_5570");
    Operation_IFC mod_5571_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5571 <- mkDebugOperation(mod_5571_inner, "mod_5571");
    Operation_IFC mod_5572_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5572 <- mkDebugOperation(mod_5572_inner, "mod_5572");
    Operation_IFC mod_5573_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5573 <- mkDebugOperation(mod_5573_inner, "mod_5573");
    Operation_IFC mod_5574_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5574 <- mkDebugOperation(mod_5574_inner, "mod_5574");
    Operation_IFC mod_5575_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5575 <- mkDebugOperation(mod_5575_inner, "mod_5575");
    Operation_IFC mod_5576_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5576 <- mkDebugOperation(mod_5576_inner, "mod_5576");
    Operation_IFC mod_5577_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5577 <- mkDebugOperation(mod_5577_inner, "mod_5577");
    Operation_IFC mod_5578_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5578 <- mkDebugOperation(mod_5578_inner, "mod_5578");
    Operation_IFC mod_5579_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5579 <- mkDebugOperation(mod_5579_inner, "mod_5579");
    Operation_IFC mod_5580_inner <- mkFlatten(1);
    Operation_IFC mod_5580 <- mkDebugOperation(mod_5580_inner, "mod_5580");
    Operation_IFC mod_5581_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5581 <- mkDebugOperation(mod_5581_inner, "mod_5581");
    Operation_IFC mod_5582_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5582 <- mkDebugOperation(mod_5582_inner, "mod_5582");
    Operation_IFC mod_5583_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5583 <- mkDebugOperation(mod_5583_inner, "mod_5583");
    Operation_IFC mod_5584_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5584 <- mkDebugOperation(mod_5584_inner, "mod_5584");
    Operation_IFC mod_5585_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5585 <- mkDebugOperation(mod_5585_inner, "mod_5585");
    Operation_IFC mod_5586_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5586 <- mkDebugOperation(mod_5586_inner, "mod_5586");
    Operation_IFC mod_5587_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5587 <- mkDebugOperation(mod_5587_inner, "mod_5587");
    Operation_IFC mod_5588_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5588 <- mkDebugOperation(mod_5588_inner, "mod_5588");
    Operation_IFC mod_5589_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5589 <- mkDebugOperation(mod_5589_inner, "mod_5589");
    Operation_IFC mod_5590_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5590 <- mkDebugOperation(mod_5590_inner, "mod_5590");
    Operation_IFC mod_5591_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5591 <- mkDebugOperation(mod_5591_inner, "mod_5591");
    Operation_IFC mod_5592_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5592 <- mkDebugOperation(mod_5592_inner, "mod_5592");
    Operation_IFC mod_5593_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5593 <- mkDebugOperation(mod_5593_inner, "mod_5593");
    Operation_IFC mod_5594_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5594 <- mkDebugOperation(mod_5594_inner, "mod_5594");
    Operation_IFC mod_5595_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5595 <- mkDebugOperation(mod_5595_inner, "mod_5595");
    Operation_IFC mod_5596_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5596 <- mkDebugOperation(mod_5596_inner, "mod_5596");
    Operation_IFC mod_5597_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5597 <- mkDebugOperation(mod_5597_inner, "mod_5597");
    Operation_IFC mod_5598_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5598 <- mkDebugOperation(mod_5598_inner, "mod_5598");
    Operation_IFC mod_5599_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5599 <- mkDebugOperation(mod_5599_inner, "mod_5599");
    Partition_IFC#(128) mod_5600_inner <- mkPartition(0, 128);
    Operation_IFC mod_5600 <- mkDebugOperation(mod_5600_inner.op, "mod_5600");
    Operation_IFC mod_5601_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5601 <- mkDebugOperation(mod_5601_inner, "mod_5601");
    Operation_IFC mod_5602_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5602 <- mkDebugOperation(mod_5602_inner, "mod_5602");
    Operation_IFC mod_5603_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5603 <- mkDebugOperation(mod_5603_inner, "mod_5603");
    Operation_IFC mod_5604_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5604 <- mkDebugOperation(mod_5604_inner, "mod_5604");
    Operation_IFC mod_5605_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5605 <- mkDebugOperation(mod_5605_inner, "mod_5605");
    Operation_IFC mod_5606_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5606 <- mkDebugOperation(mod_5606_inner, "mod_5606");
    Operation_IFC mod_5607_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5607 <- mkDebugOperation(mod_5607_inner, "mod_5607");
    Operation_IFC mod_5608_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5608 <- mkDebugOperation(mod_5608_inner, "mod_5608");
    Operation_IFC mod_5609_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5609 <- mkDebugOperation(mod_5609_inner, "mod_5609");
    Operation_IFC mod_5610_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5610 <- mkDebugOperation(mod_5610_inner, "mod_5610");
    Operation_IFC mod_5611_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5611 <- mkDebugOperation(mod_5611_inner, "mod_5611");
    Operation_IFC mod_5612_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5612 <- mkDebugOperation(mod_5612_inner, "mod_5612");
    Operation_IFC mod_5613_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5613 <- mkDebugOperation(mod_5613_inner, "mod_5613");
    Operation_IFC mod_5614_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5614 <- mkDebugOperation(mod_5614_inner, "mod_5614");
    Operation_IFC mod_5615_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5615 <- mkDebugOperation(mod_5615_inner, "mod_5615");
    Operation_IFC mod_5616_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5616 <- mkDebugOperation(mod_5616_inner, "mod_5616");
    Operation_IFC mod_5617_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5617 <- mkDebugOperation(mod_5617_inner, "mod_5617");
    Operation_IFC mod_5618_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5618 <- mkDebugOperation(mod_5618_inner, "mod_5618");
    Operation_IFC mod_5619_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5619 <- mkDebugOperation(mod_5619_inner, "mod_5619");
    Operation_IFC mod_5620_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5620 <- mkDebugOperation(mod_5620_inner, "mod_5620");
    Operation_IFC mod_5621_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5621 <- mkDebugOperation(mod_5621_inner, "mod_5621");
    Operation_IFC mod_5622_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5622 <- mkDebugOperation(mod_5622_inner, "mod_5622");
    Operation_IFC mod_5623_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5623 <- mkDebugOperation(mod_5623_inner, "mod_5623");
    Operation_IFC mod_5624_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5624 <- mkDebugOperation(mod_5624_inner, "mod_5624");
    Operation_IFC mod_5625_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5625 <- mkDebugOperation(mod_5625_inner, "mod_5625");
    Operation_IFC mod_5626_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5626 <- mkDebugOperation(mod_5626_inner, "mod_5626");
    Operation_IFC mod_5627_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5627 <- mkDebugOperation(mod_5627_inner, "mod_5627");
    Operation_IFC mod_5628_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5628 <- mkDebugOperation(mod_5628_inner, "mod_5628");
    Operation_IFC mod_5629_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5629 <- mkDebugOperation(mod_5629_inner, "mod_5629");
    Operation_IFC mod_5630_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5630 <- mkDebugOperation(mod_5630_inner, "mod_5630");
    Operation_IFC mod_5631_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5631 <- mkDebugOperation(mod_5631_inner, "mod_5631");
    Operation_IFC mod_5632_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5632 <- mkDebugOperation(mod_5632_inner, "mod_5632");
    Operation_IFC mod_5633_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5633 <- mkDebugOperation(mod_5633_inner, "mod_5633");
    Operation_IFC mod_5634_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5634 <- mkDebugOperation(mod_5634_inner, "mod_5634");
    Operation_IFC mod_5635_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5635 <- mkDebugOperation(mod_5635_inner, "mod_5635");
    Operation_IFC mod_5636_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5636 <- mkDebugOperation(mod_5636_inner, "mod_5636");
    Operation_IFC mod_5637_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5637 <- mkDebugOperation(mod_5637_inner, "mod_5637");
    Operation_IFC mod_5638_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5638 <- mkDebugOperation(mod_5638_inner, "mod_5638");
    Operation_IFC mod_5639_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5639 <- mkDebugOperation(mod_5639_inner, "mod_5639");
    Operation_IFC mod_5640_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5640 <- mkDebugOperation(mod_5640_inner, "mod_5640");
    Operation_IFC mod_5641_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5641 <- mkDebugOperation(mod_5641_inner, "mod_5641");
    Operation_IFC mod_5642_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5642 <- mkDebugOperation(mod_5642_inner, "mod_5642");
    Operation_IFC mod_5643_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5643 <- mkDebugOperation(mod_5643_inner, "mod_5643");
    Operation_IFC mod_5644_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5644 <- mkDebugOperation(mod_5644_inner, "mod_5644");
    Operation_IFC mod_5645_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5645 <- mkDebugOperation(mod_5645_inner, "mod_5645");
    Operation_IFC mod_5646_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5646 <- mkDebugOperation(mod_5646_inner, "mod_5646");
    Operation_IFC mod_5647_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5647 <- mkDebugOperation(mod_5647_inner, "mod_5647");
    Operation_IFC mod_5648_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_5648 <- mkDebugOperation(mod_5648_inner, "mod_5648");
    (* descending_urgency = "rule_6785, rule_6786, rule_6787, rule_6788, rule_6789, rule_6790, rule_6791, rule_6792, rule_6793, rule_6794, rule_6795, rule_6796, rule_6797, rule_6798, rule_6799, rule_6800, rule_6801, rule_6802, rule_6803, rule_6804, rule_6805, rule_6806, rule_6807, rule_6808, rule_6809, rule_6810, rule_6811, rule_6812, rule_6813, rule_6814, rule_6815, rule_6816, rule_6817, rule_6818, rule_6819, rule_6820, rule_6821, rule_6822, rule_6823, rule_6824, rule_6825, rule_6826, rule_6827, rule_6828, rule_6829, rule_6830, rule_6831, rule_6832, rule_6833, rule_6834, rule_6835, rule_6836, rule_6837, rule_6838, rule_6839, rule_6840, rule_6841, rule_6842, rule_6843, rule_6844, rule_6845, rule_6846, rule_6847, rule_6848, rule_6849, rule_6850, rule_6851, rule_6852, rule_6853, rule_6854, rule_6855, rule_6856, rule_6857, rule_6858, rule_6859, rule_6860, rule_6861, rule_6862, rule_6863, rule_6864, rule_6865, rule_6866, rule_6867, rule_6868, rule_6869, rule_6870, rule_6871, rule_6872, rule_6873, rule_6874, rule_6875, rule_6876, rule_6877, rule_6878, rule_6879, rule_6880, rule_6881, rule_6882, rule_6883, rule_6884, rule_6885, rule_6886, rule_6887, rule_6888, rule_6889, rule_6890, rule_6891, rule_6892, rule_6893, rule_6894, rule_6895, rule_6896, rule_6897, rule_6898, rule_6899, rule_6900, rule_6901, rule_6902, rule_6903, rule_6904, rule_6905, rule_6906, rule_6907, rule_6908, rule_6909, rule_6910, rule_6911, rule_6912, rule_6913, rule_6914, rule_6915, rule_6916, rule_6917, rule_6918, rule_6919, rule_6920, rule_6921, rule_6922, rule_6923, rule_6924, rule_6925, rule_6926, rule_6927, rule_6928, rule_6929, rule_6930, rule_6931, rule_6932, rule_6933, rule_6934, rule_6935, rule_6936, rule_6937, rule_6938, rule_6939, rule_6940, rule_6941, rule_6942, rule_6943, rule_6944, rule_6945, rule_6946, rule_6947, rule_6948, rule_6949, rule_6950, rule_6951, rule_6952, rule_6953, rule_6954, rule_6955, rule_6956, rule_6957, rule_6958, rule_6959, rule_6960, rule_6961, rule_6962, rule_6963, rule_6964, rule_6965, rule_6966, rule_6967, rule_6968, rule_6969, rule_6970, rule_6971, rule_6972, rule_6973, rule_6974, rule_6975, rule_6976, rule_6977, rule_6978, rule_6979, rule_6980, rule_6981, rule_6982, rule_6983, rule_6984, rule_6985, rule_6986, rule_6987, rule_6988, rule_6989, rule_6990, rule_6991, rule_6992, rule_6993, rule_6994, rule_6995, rule_6996, rule_6997, rule_6998, rule_6999, rule_7000, rule_7001, rule_7002, rule_7003, rule_7004, rule_7005, rule_7006, rule_7007, rule_7008, rule_7009, rule_7010, rule_7011, rule_7012, rule_7013, rule_7014, rule_7015, rule_7016, rule_7017, rule_7018, rule_7019, rule_7020, rule_7021, rule_7022, rule_7023, rule_7024, rule_7025, rule_7026, rule_7027, rule_7028, rule_7029, rule_7030, rule_7031, rule_7032, rule_7033, rule_7034, rule_7035, rule_7036, rule_7037, rule_7038, rule_7039, rule_7040, rule_7041, rule_7042, rule_7043, rule_7044, rule_7045, rule_7046, rule_7047, rule_7048, rule_7049, rule_7050, rule_7051, rule_7052, rule_7053, rule_7054, rule_7055, rule_7056, rule_7057, rule_7058, rule_7059, rule_7060, rule_7061, rule_7062, rule_7063, rule_7064, rule_7065, rule_7066, rule_7067, rule_7068, rule_7069, rule_7070, rule_7071, rule_7072, rule_7073, rule_7074, rule_7075, rule_7076, rule_7077, rule_7078, rule_7079, rule_7080, rule_7081, rule_7082, rule_7083, rule_7084, rule_7085, rule_7086, rule_7087, rule_7088, rule_7089, rule_7090, rule_7091, rule_7092, rule_7093, rule_7094, rule_7095, rule_7096, rule_7097, rule_7098, rule_7099, rule_7100, rule_7101, rule_7102, rule_7103, rule_7104, rule_7105, rule_7106, rule_7107, rule_7108, rule_7109, rule_7110, rule_7111, rule_7112, rule_7113, rule_7114, rule_7115, rule_7116, rule_7117, rule_7118, rule_7119, rule_7120, rule_7121, rule_7122, rule_7123, rule_7124, rule_7125, rule_7126, rule_7127, rule_7128, rule_7129, rule_7130, rule_7131, rule_7132, rule_7133, rule_7134, rule_7135, rule_7136, rule_7137, rule_7138, rule_7139, rule_7140, rule_7141, rule_7142, rule_7143, rule_7144, rule_7145, rule_7146, rule_7147, rule_7148, rule_7149, rule_7150, rule_7151, rule_7152, rule_7153, rule_7154, rule_7155, rule_7156, rule_7157, rule_7158, rule_7159, rule_7160, rule_7161, rule_7162, rule_7163, rule_7164, rule_7165, rule_7166, rule_7167, rule_7168, rule_7169, rule_7170, rule_7171, rule_7172, rule_7173, rule_7174, rule_7175, rule_7176, rule_7177, rule_7178, rule_7179, rule_7180, rule_7181, rule_7182, rule_7183, rule_7184, rule_7185, rule_7186, rule_7187, rule_7188, rule_7189, rule_7190, rule_7191, rule_7192, rule_7193, rule_7194, rule_7195, rule_7196, rule_7197, rule_7198, rule_7199, rule_7200, rule_7201, rule_7202, rule_7203, rule_7204, rule_7205, rule_7206, rule_7207, rule_7208, rule_7209, rule_7210, rule_7211, rule_7212, rule_7213, rule_7214, rule_7215, rule_7216, rule_7217, rule_7218, rule_7219, rule_7220, rule_7221, rule_7222, rule_7223, rule_7224, rule_7225, rule_7226, rule_7227, rule_7228, rule_7229, rule_7230, rule_7231, rule_7232, rule_7233, rule_7234, rule_7235, rule_7236, rule_7237, rule_7238, rule_7239, rule_7240, rule_7241, rule_7242, rule_7243, rule_7244, rule_7245, rule_7246, rule_7247, rule_7248, rule_7249, rule_7250, rule_7251, rule_7252, rule_7253, rule_7254, rule_7255, rule_7256, rule_7257, rule_7258, rule_7259, rule_7260, rule_7261, rule_7262, rule_7263, rule_7264, rule_7265, rule_7266, rule_7267, rule_7268, rule_7269, rule_7270, rule_7271, rule_7272, rule_7273, rule_7274, rule_7275, rule_7276, rule_7277, rule_7278, rule_7279, rule_7280, rule_7281, rule_7282, rule_7283, rule_7284, rule_7285, rule_7286, rule_7287, rule_7288, rule_7289, rule_7290, rule_7291, rule_7292, rule_7293, rule_7294, rule_7295, rule_7296, rule_7297, rule_7298, rule_7299, rule_7300, rule_7301, rule_7302, rule_7303, rule_7304, rule_7305, rule_7306, rule_7307, rule_7308, rule_7309, rule_7310, rule_7311, rule_7312, rule_7313, rule_7314, rule_7315, rule_7316, rule_7317, rule_7318, rule_7319, rule_7320, rule_7321, rule_7322, rule_7323, rule_7324, rule_7325, rule_7326, rule_7327, rule_7328, rule_7329, rule_7330, rule_7331, rule_7332, rule_7333, rule_7334, rule_7335, rule_7336, rule_7337, rule_7338, rule_7339, rule_7340, rule_7341, rule_7342, rule_7343, rule_7344, rule_7345, rule_7346, rule_7347, rule_7348, rule_7349, rule_7350, rule_7351, rule_7352, rule_7353, rule_7354, rule_7355, rule_7356, rule_7357, rule_7358, rule_7359, rule_7360, rule_7361, rule_7362, rule_7363, rule_7364, rule_7365, rule_7366, rule_7367, rule_7368, rule_7369, rule_7370, rule_7371, rule_7372, rule_7373, rule_7374, rule_7375, rule_7376, rule_7377, rule_7378, rule_7379, rule_7380, rule_7381, rule_7382, rule_7383, rule_7384, rule_7385, rule_7386, rule_7387, rule_7388, rule_7389, rule_7390, rule_7391, rule_7392, rule_7393, rule_7394, rule_7395, rule_7396, rule_7397, rule_7398, rule_7399, rule_7400, rule_7401, rule_7402, rule_7403, rule_7404, rule_7405, rule_7406, rule_7407, rule_7408, rule_7409, rule_7410, rule_7411, rule_7412, rule_7413, rule_7414, rule_7415, rule_7416, rule_7417, rule_7418, rule_7419, rule_7420, rule_7421, rule_7422, rule_7423, rule_7424, rule_7425, rule_7426, rule_7427, rule_7428, rule_7429, rule_7430, rule_7431, rule_7432, rule_7433, rule_7434, rule_7435, rule_7436, rule_7437, rule_7438, rule_7439, rule_7440, rule_7441, rule_7442, rule_7443, rule_7444, rule_7445, rule_7446, rule_7447, rule_7448, rule_7449, rule_7450, rule_7451, rule_7452, rule_7453, rule_7454, rule_7455, rule_7456, rule_7457, rule_7458, rule_7459, rule_7460, rule_7461, rule_7462, rule_7463, rule_7464, rule_7465, rule_7466, rule_7467, rule_7468, rule_7469, rule_7470, rule_7471, rule_7472, rule_7473, rule_7474, rule_7475, rule_7476, rule_7477, rule_7478, rule_7479, rule_7480, rule_7481, rule_7482, rule_7483, rule_7484, rule_7485, rule_7486, rule_7487, rule_7488, rule_7489, rule_7490, rule_7491, rule_7492, rule_7493, rule_7494, rule_7495, rule_7496, rule_7497, rule_7498, rule_7499, rule_7500, rule_7501, rule_7502, rule_7503, rule_7504, rule_7505, rule_7506, rule_7507, rule_7508, rule_7509, rule_7510, rule_7511, rule_7512, rule_7513, rule_7514, rule_7515, rule_7516, rule_7517, rule_7518, rule_7519, rule_7520, rule_7521, rule_7522, rule_7523, rule_7524, rule_7525, rule_7526, rule_7527, rule_7528, rule_7529, rule_7530, rule_7531, rule_7532, rule_7533, rule_7534, rule_7535, rule_7536, rule_7537, rule_7538, rule_7539, rule_7540, rule_7541, rule_7542, rule_7543, rule_7544, rule_7545, rule_7546, rule_7547, rule_7548, rule_7549, rule_7550, rule_7551, rule_7552, rule_7553, rule_7554, rule_7555, rule_7556, rule_7557, rule_7558, rule_7559, rule_7560, rule_7561, rule_7562, rule_7563, rule_7564, rule_7565, rule_7566, rule_7567, rule_7568, rule_7569, rule_7570, rule_7571, rule_7572, rule_7573, rule_7574, rule_7575, rule_7576, rule_7577, rule_7578, rule_7579, rule_7580, rule_7581, rule_7582, rule_7583, rule_7584, rule_7585, rule_7586, rule_7587, rule_7588, rule_7589, rule_7590, rule_7591, rule_7592, rule_7593, rule_7594, rule_7595, rule_7596, rule_7597, rule_7598, rule_7599, rule_7600, rule_7601, rule_7602, rule_7603, rule_7604, rule_7605, rule_7606, rule_7607, rule_7608, rule_7609, rule_7610, rule_7611, rule_7612, rule_7613, rule_7614, rule_7615, rule_7616, rule_7617, rule_7618, rule_7619, rule_7620, rule_7621, rule_7622, rule_7623, rule_7624, rule_7625, rule_7626, rule_7627, rule_7628, rule_7629, rule_7630, rule_7631, rule_7632, rule_7633, rule_7634, rule_7635, rule_7636, rule_7637, rule_7638, rule_7639, rule_7640, rule_7641, rule_7642, rule_7643, rule_7644, rule_7645, rule_7646, rule_7647, rule_7648, rule_7649, rule_7650, rule_7651, rule_7652, rule_7653, rule_7654, rule_7655, rule_7656, rule_7657, rule_7658, rule_7659, rule_7660, rule_7661, rule_7662, rule_7663, rule_7664, rule_7665, rule_7666, rule_7667, rule_7668, rule_7669, rule_7670, rule_7671, rule_7672, rule_7673, rule_7674, rule_7675, rule_7676, rule_7677, rule_7678, rule_7679, rule_7680, rule_7681, rule_7682, rule_7683, rule_7684, rule_7685, rule_7686, rule_7687, rule_7688, rule_7689, rule_7690, rule_7691, rule_7692, rule_7693, rule_7694, rule_7695, rule_7696, rule_7697, rule_7698, rule_7699, rule_7700, rule_7701, rule_7702, rule_7703, rule_7704, rule_7705, rule_7706, rule_7707, rule_7708, rule_7709, rule_7710, rule_7711, rule_7712, rule_7713, rule_7714, rule_7715, rule_7716, rule_7717, rule_7718, rule_7719, rule_7720, rule_7721, rule_7722, rule_7723, rule_7724, rule_7725, rule_7726, rule_7727, rule_7728, rule_7729, rule_7730, rule_7731, rule_7732, rule_7733, rule_7734, rule_7735, rule_7736, rule_7737, rule_7738, rule_7739, rule_7740, rule_7741, rule_7742, rule_7743, rule_7744, rule_7745, rule_7746, rule_7747, rule_7748, rule_7749, rule_7750, rule_7751, rule_7752, rule_7753, rule_7754, rule_7755, rule_7756, rule_7757, rule_7758, rule_7759, rule_7760, rule_7761, rule_7762, rule_7763, rule_7764, rule_7765, rule_7766, rule_7767, rule_7768, rule_7769, rule_7770, rule_7771, rule_7772, rule_7773, rule_7774, rule_7775, rule_7776, rule_7777, rule_7778, rule_7779, rule_7780, rule_7781, rule_7782, rule_7783, rule_7784, rule_7785, rule_7786, rule_7787, rule_7788, rule_7789, rule_7790, rule_7791, rule_7792, rule_7793, rule_7794, rule_7795, rule_7796, rule_7797, rule_7798, rule_7799, rule_7800, rule_7801, rule_7802, rule_7803, rule_7804, rule_7805, rule_7806, rule_7807, rule_7808, rule_7809, rule_7810, rule_7811, rule_7812, rule_7813, rule_7814, rule_7815, rule_7816, rule_7817, rule_7818, rule_7819, rule_7820, rule_7821, rule_7822, rule_7823, rule_7824, rule_7825, rule_7826, rule_7827, rule_7828, rule_7829, rule_7830, rule_7831, rule_7832, rule_7833, rule_7834, rule_7835, rule_7836, rule_7837, rule_7838, rule_7839, rule_7840, rule_7841, rule_7842, rule_7843, rule_7844, rule_7845, rule_7846, rule_7847, rule_7848, rule_7849, rule_7850, rule_7851, rule_7852, rule_7853, rule_7854, rule_7855, rule_7856, rule_7857, rule_7858, rule_7859, rule_7860, rule_7861, rule_7862, rule_7863, rule_7864, rule_7865, rule_7866, rule_7867, rule_7868, rule_7869, rule_7870, rule_7871, rule_7872, rule_7873, rule_7874, rule_7875, rule_7876, rule_7877, rule_7878, rule_7879, rule_7880, rule_7881, rule_7882, rule_7883, rule_7884, rule_7885, rule_7886, rule_7887, rule_7888, rule_7889, rule_7890, rule_7891, rule_7892, rule_7893, rule_7894, rule_7895, rule_7896, rule_7897, rule_7898, rule_7899, rule_7900, rule_7901, rule_7902, rule_7903, rule_7904, rule_7905, rule_7906, rule_7907, rule_7908, rule_7909, rule_7910, rule_7911, rule_7912, rule_7913, rule_7914, rule_7915, rule_7916, rule_7917, rule_7918, rule_7919, rule_7920, rule_7921, rule_7922, rule_7923, rule_7924, rule_7925, rule_7926, rule_7927, rule_7928, rule_7929, rule_7930, rule_7931, rule_7932, rule_7933, rule_7934, rule_7935, rule_7936, rule_7937, rule_7938, rule_7939, rule_7940, rule_7941, rule_7942, rule_7943, rule_7944, rule_7945, rule_7946, rule_7947, rule_7948, rule_7949, rule_7950, rule_7951, rule_7952" *)
    (* execution_order = "rule_6785, rule_6786, rule_6787, rule_6788, rule_6789, rule_6790, rule_6791, rule_6792, rule_6793, rule_6794, rule_6795, rule_6796, rule_6797, rule_6798, rule_6799, rule_6800, rule_6801, rule_6802, rule_6803, rule_6804, rule_6805, rule_6806, rule_6807, rule_6808, rule_6809, rule_6810, rule_6811, rule_6812, rule_6813, rule_6814, rule_6815, rule_6816, rule_6817, rule_6818, rule_6819, rule_6820, rule_6821, rule_6822, rule_6823, rule_6824, rule_6825, rule_6826, rule_6827, rule_6828, rule_6829, rule_6830, rule_6831, rule_6832, rule_6833, rule_6834, rule_6835, rule_6836, rule_6837, rule_6838, rule_6839, rule_6840, rule_6841, rule_6842, rule_6843, rule_6844, rule_6845, rule_6846, rule_6847, rule_6848, rule_6849, rule_6850, rule_6851, rule_6852, rule_6853, rule_6854, rule_6855, rule_6856, rule_6857, rule_6858, rule_6859, rule_6860, rule_6861, rule_6862, rule_6863, rule_6864, rule_6865, rule_6866, rule_6867, rule_6868, rule_6869, rule_6870, rule_6871, rule_6872, rule_6873, rule_6874, rule_6875, rule_6876, rule_6877, rule_6878, rule_6879, rule_6880, rule_6881, rule_6882, rule_6883, rule_6884, rule_6885, rule_6886, rule_6887, rule_6888, rule_6889, rule_6890, rule_6891, rule_6892, rule_6893, rule_6894, rule_6895, rule_6896, rule_6897, rule_6898, rule_6899, rule_6900, rule_6901, rule_6902, rule_6903, rule_6904, rule_6905, rule_6906, rule_6907, rule_6908, rule_6909, rule_6910, rule_6911, rule_6912, rule_6913, rule_6914, rule_6915, rule_6916, rule_6917, rule_6918, rule_6919, rule_6920, rule_6921, rule_6922, rule_6923, rule_6924, rule_6925, rule_6926, rule_6927, rule_6928, rule_6929, rule_6930, rule_6931, rule_6932, rule_6933, rule_6934, rule_6935, rule_6936, rule_6937, rule_6938, rule_6939, rule_6940, rule_6941, rule_6942, rule_6943, rule_6944, rule_6945, rule_6946, rule_6947, rule_6948, rule_6949, rule_6950, rule_6951, rule_6952, rule_6953, rule_6954, rule_6955, rule_6956, rule_6957, rule_6958, rule_6959, rule_6960, rule_6961, rule_6962, rule_6963, rule_6964, rule_6965, rule_6966, rule_6967, rule_6968, rule_6969, rule_6970, rule_6971, rule_6972, rule_6973, rule_6974, rule_6975, rule_6976, rule_6977, rule_6978, rule_6979, rule_6980, rule_6981, rule_6982, rule_6983, rule_6984, rule_6985, rule_6986, rule_6987, rule_6988, rule_6989, rule_6990, rule_6991, rule_6992, rule_6993, rule_6994, rule_6995, rule_6996, rule_6997, rule_6998, rule_6999, rule_7000, rule_7001, rule_7002, rule_7003, rule_7004, rule_7005, rule_7006, rule_7007, rule_7008, rule_7009, rule_7010, rule_7011, rule_7012, rule_7013, rule_7014, rule_7015, rule_7016, rule_7017, rule_7018, rule_7019, rule_7020, rule_7021, rule_7022, rule_7023, rule_7024, rule_7025, rule_7026, rule_7027, rule_7028, rule_7029, rule_7030, rule_7031, rule_7032, rule_7033, rule_7034, rule_7035, rule_7036, rule_7037, rule_7038, rule_7039, rule_7040, rule_7041, rule_7042, rule_7043, rule_7044, rule_7045, rule_7046, rule_7047, rule_7048, rule_7049, rule_7050, rule_7051, rule_7052, rule_7053, rule_7054, rule_7055, rule_7056, rule_7057, rule_7058, rule_7059, rule_7060, rule_7061, rule_7062, rule_7063, rule_7064, rule_7065, rule_7066, rule_7067, rule_7068, rule_7069, rule_7070, rule_7071, rule_7072, rule_7073, rule_7074, rule_7075, rule_7076, rule_7077, rule_7078, rule_7079, rule_7080, rule_7081, rule_7082, rule_7083, rule_7084, rule_7085, rule_7086, rule_7087, rule_7088, rule_7089, rule_7090, rule_7091, rule_7092, rule_7093, rule_7094, rule_7095, rule_7096, rule_7097, rule_7098, rule_7099, rule_7100, rule_7101, rule_7102, rule_7103, rule_7104, rule_7105, rule_7106, rule_7107, rule_7108, rule_7109, rule_7110, rule_7111, rule_7112, rule_7113, rule_7114, rule_7115, rule_7116, rule_7117, rule_7118, rule_7119, rule_7120, rule_7121, rule_7122, rule_7123, rule_7124, rule_7125, rule_7126, rule_7127, rule_7128, rule_7129, rule_7130, rule_7131, rule_7132, rule_7133, rule_7134, rule_7135, rule_7136, rule_7137, rule_7138, rule_7139, rule_7140, rule_7141, rule_7142, rule_7143, rule_7144, rule_7145, rule_7146, rule_7147, rule_7148, rule_7149, rule_7150, rule_7151, rule_7152, rule_7153, rule_7154, rule_7155, rule_7156, rule_7157, rule_7158, rule_7159, rule_7160, rule_7161, rule_7162, rule_7163, rule_7164, rule_7165, rule_7166, rule_7167, rule_7168, rule_7169, rule_7170, rule_7171, rule_7172, rule_7173, rule_7174, rule_7175, rule_7176, rule_7177, rule_7178, rule_7179, rule_7180, rule_7181, rule_7182, rule_7183, rule_7184, rule_7185, rule_7186, rule_7187, rule_7188, rule_7189, rule_7190, rule_7191, rule_7192, rule_7193, rule_7194, rule_7195, rule_7196, rule_7197, rule_7198, rule_7199, rule_7200, rule_7201, rule_7202, rule_7203, rule_7204, rule_7205, rule_7206, rule_7207, rule_7208, rule_7209, rule_7210, rule_7211, rule_7212, rule_7213, rule_7214, rule_7215, rule_7216, rule_7217, rule_7218, rule_7219, rule_7220, rule_7221, rule_7222, rule_7223, rule_7224, rule_7225, rule_7226, rule_7227, rule_7228, rule_7229, rule_7230, rule_7231, rule_7232, rule_7233, rule_7234, rule_7235, rule_7236, rule_7237, rule_7238, rule_7239, rule_7240, rule_7241, rule_7242, rule_7243, rule_7244, rule_7245, rule_7246, rule_7247, rule_7248, rule_7249, rule_7250, rule_7251, rule_7252, rule_7253, rule_7254, rule_7255, rule_7256, rule_7257, rule_7258, rule_7259, rule_7260, rule_7261, rule_7262, rule_7263, rule_7264, rule_7265, rule_7266, rule_7267, rule_7268, rule_7269, rule_7270, rule_7271, rule_7272, rule_7273, rule_7274, rule_7275, rule_7276, rule_7277, rule_7278, rule_7279, rule_7280, rule_7281, rule_7282, rule_7283, rule_7284, rule_7285, rule_7286, rule_7287, rule_7288, rule_7289, rule_7290, rule_7291, rule_7292, rule_7293, rule_7294, rule_7295, rule_7296, rule_7297, rule_7298, rule_7299, rule_7300, rule_7301, rule_7302, rule_7303, rule_7304, rule_7305, rule_7306, rule_7307, rule_7308, rule_7309, rule_7310, rule_7311, rule_7312, rule_7313, rule_7314, rule_7315, rule_7316, rule_7317, rule_7318, rule_7319, rule_7320, rule_7321, rule_7322, rule_7323, rule_7324, rule_7325, rule_7326, rule_7327, rule_7328, rule_7329, rule_7330, rule_7331, rule_7332, rule_7333, rule_7334, rule_7335, rule_7336, rule_7337, rule_7338, rule_7339, rule_7340, rule_7341, rule_7342, rule_7343, rule_7344, rule_7345, rule_7346, rule_7347, rule_7348, rule_7349, rule_7350, rule_7351, rule_7352, rule_7353, rule_7354, rule_7355, rule_7356, rule_7357, rule_7358, rule_7359, rule_7360, rule_7361, rule_7362, rule_7363, rule_7364, rule_7365, rule_7366, rule_7367, rule_7368, rule_7369, rule_7370, rule_7371, rule_7372, rule_7373, rule_7374, rule_7375, rule_7376, rule_7377, rule_7378, rule_7379, rule_7380, rule_7381, rule_7382, rule_7383, rule_7384, rule_7385, rule_7386, rule_7387, rule_7388, rule_7389, rule_7390, rule_7391, rule_7392, rule_7393, rule_7394, rule_7395, rule_7396, rule_7397, rule_7398, rule_7399, rule_7400, rule_7401, rule_7402, rule_7403, rule_7404, rule_7405, rule_7406, rule_7407, rule_7408, rule_7409, rule_7410, rule_7411, rule_7412, rule_7413, rule_7414, rule_7415, rule_7416, rule_7417, rule_7418, rule_7419, rule_7420, rule_7421, rule_7422, rule_7423, rule_7424, rule_7425, rule_7426, rule_7427, rule_7428, rule_7429, rule_7430, rule_7431, rule_7432, rule_7433, rule_7434, rule_7435, rule_7436, rule_7437, rule_7438, rule_7439, rule_7440, rule_7441, rule_7442, rule_7443, rule_7444, rule_7445, rule_7446, rule_7447, rule_7448, rule_7449, rule_7450, rule_7451, rule_7452, rule_7453, rule_7454, rule_7455, rule_7456, rule_7457, rule_7458, rule_7459, rule_7460, rule_7461, rule_7462, rule_7463, rule_7464, rule_7465, rule_7466, rule_7467, rule_7468, rule_7469, rule_7470, rule_7471, rule_7472, rule_7473, rule_7474, rule_7475, rule_7476, rule_7477, rule_7478, rule_7479, rule_7480, rule_7481, rule_7482, rule_7483, rule_7484, rule_7485, rule_7486, rule_7487, rule_7488, rule_7489, rule_7490, rule_7491, rule_7492, rule_7493, rule_7494, rule_7495, rule_7496, rule_7497, rule_7498, rule_7499, rule_7500, rule_7501, rule_7502, rule_7503, rule_7504, rule_7505, rule_7506, rule_7507, rule_7508, rule_7509, rule_7510, rule_7511, rule_7512, rule_7513, rule_7514, rule_7515, rule_7516, rule_7517, rule_7518, rule_7519, rule_7520, rule_7521, rule_7522, rule_7523, rule_7524, rule_7525, rule_7526, rule_7527, rule_7528, rule_7529, rule_7530, rule_7531, rule_7532, rule_7533, rule_7534, rule_7535, rule_7536, rule_7537, rule_7538, rule_7539, rule_7540, rule_7541, rule_7542, rule_7543, rule_7544, rule_7545, rule_7546, rule_7547, rule_7548, rule_7549, rule_7550, rule_7551, rule_7552, rule_7553, rule_7554, rule_7555, rule_7556, rule_7557, rule_7558, rule_7559, rule_7560, rule_7561, rule_7562, rule_7563, rule_7564, rule_7565, rule_7566, rule_7567, rule_7568, rule_7569, rule_7570, rule_7571, rule_7572, rule_7573, rule_7574, rule_7575, rule_7576, rule_7577, rule_7578, rule_7579, rule_7580, rule_7581, rule_7582, rule_7583, rule_7584, rule_7585, rule_7586, rule_7587, rule_7588, rule_7589, rule_7590, rule_7591, rule_7592, rule_7593, rule_7594, rule_7595, rule_7596, rule_7597, rule_7598, rule_7599, rule_7600, rule_7601, rule_7602, rule_7603, rule_7604, rule_7605, rule_7606, rule_7607, rule_7608, rule_7609, rule_7610, rule_7611, rule_7612, rule_7613, rule_7614, rule_7615, rule_7616, rule_7617, rule_7618, rule_7619, rule_7620, rule_7621, rule_7622, rule_7623, rule_7624, rule_7625, rule_7626, rule_7627, rule_7628, rule_7629, rule_7630, rule_7631, rule_7632, rule_7633, rule_7634, rule_7635, rule_7636, rule_7637, rule_7638, rule_7639, rule_7640, rule_7641, rule_7642, rule_7643, rule_7644, rule_7645, rule_7646, rule_7647, rule_7648, rule_7649, rule_7650, rule_7651, rule_7652, rule_7653, rule_7654, rule_7655, rule_7656, rule_7657, rule_7658, rule_7659, rule_7660, rule_7661, rule_7662, rule_7663, rule_7664, rule_7665, rule_7666, rule_7667, rule_7668, rule_7669, rule_7670, rule_7671, rule_7672, rule_7673, rule_7674, rule_7675, rule_7676, rule_7677, rule_7678, rule_7679, rule_7680, rule_7681, rule_7682, rule_7683, rule_7684, rule_7685, rule_7686, rule_7687, rule_7688, rule_7689, rule_7690, rule_7691, rule_7692, rule_7693, rule_7694, rule_7695, rule_7696, rule_7697, rule_7698, rule_7699, rule_7700, rule_7701, rule_7702, rule_7703, rule_7704, rule_7705, rule_7706, rule_7707, rule_7708, rule_7709, rule_7710, rule_7711, rule_7712, rule_7713, rule_7714, rule_7715, rule_7716, rule_7717, rule_7718, rule_7719, rule_7720, rule_7721, rule_7722, rule_7723, rule_7724, rule_7725, rule_7726, rule_7727, rule_7728, rule_7729, rule_7730, rule_7731, rule_7732, rule_7733, rule_7734, rule_7735, rule_7736, rule_7737, rule_7738, rule_7739, rule_7740, rule_7741, rule_7742, rule_7743, rule_7744, rule_7745, rule_7746, rule_7747, rule_7748, rule_7749, rule_7750, rule_7751, rule_7752, rule_7753, rule_7754, rule_7755, rule_7756, rule_7757, rule_7758, rule_7759, rule_7760, rule_7761, rule_7762, rule_7763, rule_7764, rule_7765, rule_7766, rule_7767, rule_7768, rule_7769, rule_7770, rule_7771, rule_7772, rule_7773, rule_7774, rule_7775, rule_7776, rule_7777, rule_7778, rule_7779, rule_7780, rule_7781, rule_7782, rule_7783, rule_7784, rule_7785, rule_7786, rule_7787, rule_7788, rule_7789, rule_7790, rule_7791, rule_7792, rule_7793, rule_7794, rule_7795, rule_7796, rule_7797, rule_7798, rule_7799, rule_7800, rule_7801, rule_7802, rule_7803, rule_7804, rule_7805, rule_7806, rule_7807, rule_7808, rule_7809, rule_7810, rule_7811, rule_7812, rule_7813, rule_7814, rule_7815, rule_7816, rule_7817, rule_7818, rule_7819, rule_7820, rule_7821, rule_7822, rule_7823, rule_7824, rule_7825, rule_7826, rule_7827, rule_7828, rule_7829, rule_7830, rule_7831, rule_7832, rule_7833, rule_7834, rule_7835, rule_7836, rule_7837, rule_7838, rule_7839, rule_7840, rule_7841, rule_7842, rule_7843, rule_7844, rule_7845, rule_7846, rule_7847, rule_7848, rule_7849, rule_7850, rule_7851, rule_7852, rule_7853, rule_7854, rule_7855, rule_7856, rule_7857, rule_7858, rule_7859, rule_7860, rule_7861, rule_7862, rule_7863, rule_7864, rule_7865, rule_7866, rule_7867, rule_7868, rule_7869, rule_7870, rule_7871, rule_7872, rule_7873, rule_7874, rule_7875, rule_7876, rule_7877, rule_7878, rule_7879, rule_7880, rule_7881, rule_7882, rule_7883, rule_7884, rule_7885, rule_7886, rule_7887, rule_7888, rule_7889, rule_7890, rule_7891, rule_7892, rule_7893, rule_7894, rule_7895, rule_7896, rule_7897, rule_7898, rule_7899, rule_7900, rule_7901, rule_7902, rule_7903, rule_7904, rule_7905, rule_7906, rule_7907, rule_7908, rule_7909, rule_7910, rule_7911, rule_7912, rule_7913, rule_7914, rule_7915, rule_7916, rule_7917, rule_7918, rule_7919, rule_7920, rule_7921, rule_7922, rule_7923, rule_7924, rule_7925, rule_7926, rule_7927, rule_7928, rule_7929, rule_7930, rule_7931, rule_7932, rule_7933, rule_7934, rule_7935, rule_7936, rule_7937, rule_7938, rule_7939, rule_7940, rule_7941, rule_7942, rule_7943, rule_7944, rule_7945, rule_7946, rule_7947, rule_7948, rule_7949, rule_7950, rule_7951, rule_7952" *)
    rule rule_6785;
        ChannelMessage t;
        t <- mod_5532.get(0);
        mod_4633.put(3, t);
    endrule
    rule rule_6786;
        ChannelMessage t;
        t <- mod_5600.get(4);
        mod_164.put(1, t);
    endrule
    rule rule_6787;
        ChannelMessage t;
        t <- mod_5451.get(0);
        mod_1025.put(2, t);
    endrule
    rule rule_6788;
        ChannelMessage t;
        t <- mod_5457.get(0);
        mod_4182.put(4, t);
    endrule
    rule rule_6789;
        ChannelMessage t;
        t <- mod_902.get(0);
        mod_5382.put(0, t);
    endrule
    rule rule_6790;
        ChannelMessage t;
        t <- mod_984.get(0);
        mod_5313.put(103, t);
    endrule
    rule rule_6791;
        ChannelMessage t;
        t <- mod_3321.get(1);
        mod_5313.put(46, t);
    endrule
    rule rule_6792;
        ChannelMessage t;
        t <- mod_5309.get(93);
        mod_3813.put(0, t);
    endrule
    rule rule_6793;
        ChannelMessage t;
        t <- mod_3608.get(3);
        mod_5401.put(0, t);
    endrule
    rule rule_6794;
        ChannelMessage t;
        t <- mod_5565.get(0);
        mod_4633.put(4, t);
    endrule
    rule rule_6795;
        ChannelMessage t;
        t <- mod_5329.get(0);
        mod_1845.put(4, t);
    endrule
    rule rule_6796;
        ChannelMessage t;
        t <- mod_5309.get(55);
        mod_2255.put(0, t);
    endrule
    rule rule_6797;
        ChannelMessage t;
        t <- mod_5402.get(0);
        mod_3690.put(4, t);
    endrule
    rule rule_6798;
        ChannelMessage t;
        t <- mod_5627.get(0);
        mod_4428.put(3, t);
    endrule
    rule rule_6799;
        ChannelMessage t;
        t <- mod_5584.get(0);
        mod_1517.put(3, t);
    endrule
    rule rule_6800;
        ChannelMessage t;
        t <- mod_5648.get(0);
        mod_2460.put(2, t);
    endrule
    rule rule_6801;
        ChannelMessage t;
        t <- mod_5326.get(1);
        mod_5372.put(1, t);
    endrule
    rule rule_6802;
        ChannelMessage t;
        t <- mod_2214.get(3);
        mod_5420.put(0, t);
    endrule
    rule rule_6803;
        ChannelMessage t;
        t <- mod_5309.get(101);
        mod_4141.put(0, t);
    endrule
    rule rule_6804;
        ChannelMessage t;
        t <- mod_1927.get(1);
        mod_5310.put(0, t);
    endrule
    rule rule_6805;
        ChannelMessage t;
        t <- mod_5390.get(0);
        mod_1230.put(4, t);
    endrule
    rule rule_6806;
        ChannelMessage t;
        t <- mod_5364.get(0);
        mod_2255.put(3, t);
    endrule
    rule rule_6807;
        ChannelMessage t;
        t <- mod_5500.get(0);
        mod_123.put(3, t);
    endrule
    rule rule_6808;
        ChannelMessage t;
        t <- mod_5309.get(107);
        mod_4387.put(0, t);
    endrule
    rule rule_6809;
        ChannelMessage t;
        t <- mod_82.get(1);
        mod_5272.put(0, t);
    endrule
    rule rule_6810;
        ChannelMessage t;
        t <- mod_4510.get(3);
        mod_5558.put(0, t);
    endrule
    rule rule_6811;
        ChannelMessage t;
        t <- mod_5600.get(116);
        mod_4756.put(1, t);
    endrule
    rule rule_6812;
        ChannelMessage t;
        t <- mod_1599.get(0);
        mod_5313.put(88, t);
    endrule
    rule rule_6813;
        ChannelMessage t;
        t <- mod_3813.get(1);
        mod_5345.put(0, t);
    endrule
    rule rule_6814;
        ChannelMessage t;
        t <- mod_5496.get(0);
        mod_3731.put(3, t);
    endrule
    rule rule_6815;
        ChannelMessage t;
        t <- mod_5309.get(62);
        mod_2542.put(0, t);
    endrule
    rule rule_6816;
        ChannelMessage t;
        t <- mod_5380.get(0);
        mod_1312.put(3, t);
    endrule
    rule rule_6817;
        ChannelMessage t;
        t <- mod_5461.get(0);
        mod_246.put(3, t);
    endrule
    rule rule_6818;
        ChannelMessage t;
        t <- mod_5309.get(118);
        mod_4838.put(0, t);
    endrule
    rule rule_6819;
        ChannelMessage t;
        t <- mod_5589.get(0);
        mod_1558.put(2, t);
    endrule
    rule rule_6820;
        ChannelMessage t;
        t <- mod_5594.get(0);
        mod_4305.put(4, t);
    endrule
    rule rule_6821;
        ChannelMessage t;
        t <- mod_5309.get(8);
        mod_328.put(0, t);
    endrule
    rule rule_6822;
        ChannelMessage t;
        t <- mod_5408.get(0);
        mod_2952.put(2, t);
    endrule
    rule rule_6823;
        ChannelMessage t;
        t <- mod_5309.get(108);
        mod_4428.put(0, t);
    endrule
    rule rule_6824;
        ChannelMessage t;
        t <- mod_5600.get(64);
        mod_2624.put(1, t);
    endrule
    rule rule_6825;
        ChannelMessage t;
        t <- mod_5600.get(88);
        mod_3608.put(1, t);
    endrule
    rule rule_6826;
        ChannelMessage t;
        t <- mod_5600.get(103);
        mod_4223.put(1, t);
    endrule
    rule rule_6827;
        ChannelMessage t;
        t <- mod_3608.get(0);
        mod_5346.put(0, t);
    endrule
    rule rule_6828;
        ChannelMessage t;
        t <- mod_5600.get(71);
        mod_2911.put(1, t);
    endrule
    rule rule_6829;
        ChannelMessage t;
        t <- mod_5587.get(0);
        mod_1722.put(2, t);
    endrule
    rule rule_6830;
        ChannelMessage t;
        t <- mod_1312.get(3);
        mod_5380.put(0, t);
    endrule
    rule rule_6831;
        ChannelMessage t;
        t <- mod_1353.get(1);
        mod_5471.put(0, t);
    endrule
    rule rule_6832;
        ChannelMessage t;
        t <- mod_5391.get(0);
        mod_4551.put(2, t);
    endrule
    rule rule_6833;
        ChannelMessage t;
        t <- mod_5600.get(87);
        mod_3567.put(1, t);
    endrule
    rule rule_6834;
        ChannelMessage t;
        t <- mod_5309.get(102);
        mod_4182.put(0, t);
    endrule
    rule rule_6835;
        ChannelMessage t;
        t <- mod_861.get(0);
        mod_5313.put(106, t);
    endrule
    rule rule_6836;
        ChannelMessage t;
        t <- mod_2337.get(1);
        mod_5313.put(70, t);
    endrule
    rule rule_6837;
        ChannelMessage t;
        t <- mod_5600.get(36);
        mod_1476.put(1, t);
    endrule
    rule rule_6838;
        ChannelMessage t;
        t <- mod_5646.get(0);
        mod_5166.put(4, t);
    endrule
    rule rule_6839;
        ChannelMessage t;
        t <- mod_5600.get(33);
        mod_1353.put(1, t);
    endrule
    rule rule_6840;
        ChannelMessage t;
        t <- mod_984.get(3);
        mod_5353.put(0, t);
    endrule
    rule rule_6841;
        ChannelMessage t;
        t <- mod_5600.get(28);
        mod_1148.put(1, t);
    endrule
    rule rule_6842;
        ChannelMessage t;
        t <- mod_1435.get(0);
        mod_5417.put(0, t);
    endrule
    rule rule_6843;
        ChannelMessage t;
        t <- mod_5309.get(115);
        mod_4715.put(0, t);
    endrule
    rule rule_6844;
        ChannelMessage t;
        t <- mod_5624.get(0);
        mod_1025.put(3, t);
    endrule
    rule rule_6845;
        ChannelMessage t;
        t <- mod_5600.get(68);
        mod_2788.put(1, t);
    endrule
    rule rule_6846;
        ChannelMessage t;
        t <- mod_4797.get(0);
        mod_5354.put(0, t);
    endrule
    rule rule_6847;
        ChannelMessage t;
        t <- mod_4838.get(0);
        mod_5313.put(9, t);
    endrule
    rule rule_6848;
        ChannelMessage t;
        t <- mod_410.get(3);
        mod_5313.put(117, t);
    endrule
    rule rule_6849;
        ChannelMessage t;
        t <- mod_5465.get(0);
        mod_1230.put(3, t);
    endrule
    rule rule_6850;
        ChannelMessage t;
        t <- mod_5600.get(80);
        mod_3280.put(1, t);
    endrule
    rule rule_6851;
        ChannelMessage t;
        t <- mod_5600.get(37);
        mod_1517.put(1, t);
    endrule
    rule rule_6852;
        ChannelMessage t;
        t <- mod_3280.get(0);
        mod_5313.put(47, t);
    endrule
    rule rule_6853;
        ChannelMessage t;
        t <- mod_3813.get(2);
        mod_5361.put(0, t);
    endrule
    rule rule_6854;
        ChannelMessage t;
        t <- mod_3567.get(0);
        mod_5606.put(0, t);
    endrule
    rule rule_6855;
        ChannelMessage t;
        t <- mod_5288.get(0);
        mod_3895.put(3, t);
    endrule
    rule rule_6856;
        ChannelMessage t;
        t <- mod_5562.get(0);
        mod_4018.put(2, t);
    endrule
    rule rule_6857;
        ChannelMessage t;
        t <- mod_5600.get(48);
        mod_1968.put(1, t);
    endrule
    rule rule_6858;
        ChannelMessage t;
        t <- mod_5426.get(0);
        mod_5523.put(0, t);
    endrule
    rule rule_6859;
        ChannelMessage t;
        t <- mod_5579.get(0);
        mod_1394.put(3, t);
    endrule
    rule rule_6860;
        ChannelMessage t;
        t <- mod_5600.get(8);
        mod_328.put(1, t);
    endrule
    rule rule_6861;
        ChannelMessage t;
        t <- mod_3321.get(0);
        mod_5641.put(0, t);
    endrule
    rule rule_6862;
        ChannelMessage t;
        t <- mod_574.get(3);
        mod_5517.put(0, t);
    endrule
    rule rule_6863;
        ChannelMessage t;
        t <- mod_5600.get(73);
        mod_2993.put(1, t);
    endrule
    rule rule_6864;
        ChannelMessage t;
        t <- mod_5600.get(110);
        mod_4510.put(1, t);
    endrule
    rule rule_6865;
        ChannelMessage t;
        t <- mod_5600.get(50);
        mod_2050.put(1, t);
    endrule
    rule rule_6866;
        ChannelMessage t;
        t <- mod_4346.get(0);
        mod_5439.put(0, t);
    endrule
    rule rule_6867;
        ChannelMessage t;
        t <- mod_5309.get(91);
        mod_3731.put(0, t);
    endrule
    rule rule_6868;
        ChannelMessage t;
        t <- mod_5419.get(0);
        mod_902.put(2, t);
    endrule
    rule rule_6869;
        ChannelMessage t;
        t <- mod_3485.get(3);
        mod_5400.put(0, t);
    endrule
    rule rule_6870;
        ChannelMessage t;
        t <- mod_3813.get(3);
        mod_5313.put(34, t);
    endrule
    rule rule_6871;
        ChannelMessage t;
        t <- mod_5125.get(0);
        mod_5313.put(2, t);
    endrule
    rule rule_6872;
        ChannelMessage t;
        t <- mod_5309.get(22);
        mod_902.put(0, t);
    endrule
    rule rule_6873;
        ChannelMessage t;
        t <- mod_3608.get(2);
        mod_5303.put(0, t);
    endrule
    rule rule_6874;
        ChannelMessage t;
        t <- mod_5309.get(63);
        mod_2583.put(0, t);
    endrule
    rule rule_6875;
        ChannelMessage t;
        t <- mod_5309.get(72);
        mod_2952.put(0, t);
    endrule
    rule rule_6876;
        ChannelMessage t;
        t <- mod_5311.get(0);
        mod_328.put(2, t);
    endrule
    rule rule_6877;
        ChannelMessage t;
        t <- mod_5492.get(0);
        mod_4633.put(2, t);
    endrule
    rule rule_6878;
        ChannelMessage t;
        t <- mod_1722.get(0);
        mod_5611.put(0, t);
    endrule
    rule rule_6879;
        ChannelMessage t;
        t <- mod_5600.get(21);
        mod_861.put(1, t);
    endrule
    rule rule_6880;
        ChannelMessage t;
        t <- mod_5341.get(0);
        mod_205.put(4, t);
    endrule
    rule rule_6881;
        ChannelMessage t;
        t <- mod_5600.get(94);
        mod_3854.put(1, t);
    endrule
    rule rule_6882;
        ChannelMessage t;
        t <- mod_5600.get(118);
        mod_4838.put(1, t);
    endrule
    rule rule_6883;
        ChannelMessage t;
        t <- mod_5608.get(0);
        mod_2829.put(4, t);
    endrule
    rule rule_6884;
        ChannelMessage t;
        t <- mod_5619.get(0);
        mod_1763.put(2, t);
    endrule
    rule rule_6885;
        ChannelMessage t;
        t <- mod_5084.get(2);
        mod_5313.put(3, t);
    endrule
    rule rule_6886;
        ChannelMessage t;
        t <- mod_5610.get(0);
        mod_492.put(4, t);
    endrule
    rule rule_6887;
        ChannelMessage t;
        t <- mod_1312.get(0);
        mod_5313.put(95, t);
    endrule
    rule rule_6888;
        ChannelMessage t;
        t <- mod_5309.get(74);
        mod_3034.put(0, t);
    endrule
    rule rule_6889;
        ChannelMessage t;
        t <- mod_5458.get(0);
        mod_4838.put(3, t);
    endrule
    rule rule_6890;
        ChannelMessage t;
        t <- mod_5166.get(2);
        mod_5313.put(1, t);
    endrule
    rule rule_6891;
        ChannelMessage t;
        t <- mod_3936.get(3);
        mod_5280.put(0, t);
    endrule
    rule rule_6892;
        ChannelMessage t;
        t <- mod_5309.get(25);
        mod_1025.put(0, t);
    endrule
    rule rule_6893;
        ChannelMessage t;
        t <- mod_820.get(2);
        mod_5405.put(0, t);
    endrule
    rule rule_6894;
        ChannelMessage t;
        t <- mod_2419.get(2);
        mod_5605.put(0, t);
    endrule
    rule rule_6895;
        ChannelMessage t;
        t <- mod_4920.get(3);
        mod_5536.put(0, t);
    endrule
    rule rule_6896;
        ChannelMessage t;
        t <- mod_5309.get(21);
        mod_861.put(0, t);
    endrule
    rule rule_6897;
        ChannelMessage t;
        t <- mod_5309.get(31);
        mod_1271.put(0, t);
    endrule
    rule rule_6898;
        ChannelMessage t;
        t <- mod_5571.get(0);
        mod_2132.put(4, t);
    endrule
    rule rule_6899;
        ChannelMessage t;
        t <- mod_5490.get(0);
        mod_943.put(4, t);
    endrule
    rule rule_6900;
        ChannelMessage t;
        t <- mod_2296.get(3);
        mod_5270.put(0, t);
    endrule
    rule rule_6901;
        ChannelMessage t;
        t <- mod_3239.get(2);
        mod_5498.put(0, t);
    endrule
    rule rule_6902;
        ChannelMessage t;
        t <- mod_5043.get(0);
        mod_5274.put(0, t);
    endrule
    rule rule_6903;
        ChannelMessage t;
        t <- mod_5600.get(29);
        mod_1189.put(1, t);
    endrule
    rule rule_6904;
        ChannelMessage t;
        t <- mod_4346.get(1);
        mod_5264.put(0, t);
    endrule
    rule rule_6905;
        ChannelMessage t;
        t <- mod_4182.get(1);
        mod_5457.put(0, t);
    endrule
    rule rule_6906;
        ChannelMessage t;
        t <- mod_5309.get(37);
        mod_1517.put(0, t);
    endrule
    rule rule_6907;
        ChannelMessage t;
        t <- mod_5298.get(0);
        mod_697.put(2, t);
    endrule
    rule rule_6908;
        ChannelMessage t;
        t <- mod_4018.get(1);
        mod_5562.put(0, t);
    endrule
    rule rule_6909;
        ChannelMessage t;
        t <- mod_5600.get(86);
        mod_3526.put(1, t);
    endrule
    rule rule_6910;
        ChannelMessage t;
        t <- mod_5309.get(75);
        mod_3075.put(0, t);
    endrule
    rule rule_6911;
        ChannelMessage t;
        t <- mod_4428.get(1);
        mod_5313.put(19, t);
    endrule
    rule rule_6912;
        ChannelMessage t;
        t <- mod_5600.get(60);
        mod_2460.put(1, t);
    endrule
    rule rule_6913;
        ChannelMessage t;
        t <- mod_5414.get(0);
        mod_1476.put(2, t);
    endrule
    rule rule_6914;
        ChannelMessage t;
        t <- mod_5527.get(0);
        mod_1640.put(4, t);
    endrule
    rule rule_6915;
        ChannelMessage t;
        t <- mod_697.get(2);
        mod_5483.put(0, t);
    endrule
    rule rule_6916;
        ChannelMessage t;
        t <- mod_4100.get(1);
        mod_5313.put(27, t);
    endrule
    rule rule_6917;
        ChannelMessage t;
        t <- mod_5600.get(102);
        mod_4182.put(1, t);
    endrule
    rule rule_6918;
        ChannelMessage t;
        t <- mod_5410.get(0);
        mod_4141.put(2, t);
    endrule
    rule rule_6919;
        ChannelMessage t;
        t <- mod_5604.get(0);
        mod_410.put(2, t);
    endrule
    rule rule_6920;
        ChannelMessage t;
        t <- mod_5352.get(0);
        mod_4100.put(2, t);
    endrule
    rule rule_6921;
        ChannelMessage t;
        t <- mod_5309.get(103);
        mod_4223.put(0, t);
    endrule
    rule rule_6922;
        ChannelMessage t;
        t <- mod_5425.get(0);
        mod_4141.put(4, t);
    endrule
    rule rule_6923;
        ChannelMessage t;
        t <- mod_1927.get(2);
        mod_5313.put(80, t);
    endrule
    rule rule_6924;
        ChannelMessage t;
        t <- mod_5600.get(3);
        mod_123.put(1, t);
    endrule
    rule rule_6925;
        ChannelMessage t;
        t <- mod_3772.get(1);
        mod_5313.put(35, t);
    endrule
    rule rule_6926;
        ChannelMessage t;
        t <- mod_5207.get(3);
        mod_5475.put(0, t);
    endrule
    rule rule_6927;
        ChannelMessage t;
        t <- mod_5375.get(0);
        mod_4674.put(2, t);
    endrule
    rule rule_6928;
        ChannelMessage t;
        t <- mod_5600.get(121);
        mod_4961.put(1, t);
    endrule
    rule rule_6929;
        ChannelMessage t;
        t <- mod_5498.get(0);
        mod_3239.put(4, t);
    endrule
    rule rule_6930;
        ChannelMessage t;
        t <- mod_5355.get(0);
        mod_3157.put(4, t);
    endrule
    rule rule_6931;
        ChannelMessage t;
        t <- mod_328.get(3);
        mod_5313.put(119, t);
    endrule
    rule rule_6932;
        ChannelMessage t;
        t <- mod_1107.get(1);
        mod_5299.put(0, t);
    endrule
    rule rule_6933;
        ChannelMessage t;
        t <- mod_5545.get(0);
        mod_2050.put(2, t);
    endrule
    rule rule_6934;
        ChannelMessage t;
        t <- mod_5309.get(29);
        mod_1189.put(0, t);
    endrule
    rule rule_6935;
        ChannelMessage t;
        t <- mod_2501.get(0);
        mod_5369.put(0, t);
    endrule
    rule rule_6936;
        ChannelMessage t;
        t <- mod_3075.get(2);
        mod_5585.put(0, t);
    endrule
    rule rule_6937;
        ChannelMessage t;
        t <- mod_5309.get(11);
        mod_451.put(0, t);
    endrule
    rule rule_6938;
        ChannelMessage t;
        t <- mod_5600.get(22);
        mod_902.put(1, t);
    endrule
    rule rule_6939;
        ChannelMessage t;
        t <- mod_5600.get(59);
        mod_2419.put(1, t);
    endrule
    rule rule_6940;
        ChannelMessage t;
        t <- mod_5455.get(0);
        mod_574.put(3, t);
    endrule
    rule rule_6941;
        ChannelMessage t;
        t <- mod_5596.get(0);
        mod_3403.put(2, t);
    endrule
    rule rule_6942;
        ChannelMessage t;
        t <- mod_1517.get(0);
        mod_5535.put(0, t);
    endrule
    rule rule_6943;
        ChannelMessage t;
        t <- mod_574.get(0);
        mod_5385.put(0, t);
    endrule
    rule rule_6944;
        ChannelMessage t;
        t <- mod_2050.get(3);
        mod_5545.put(0, t);
    endrule
    rule rule_6945;
        ChannelMessage t;
        t <- mod_4346.get(2);
        mod_5520.put(0, t);
    endrule
    rule rule_6946;
        ChannelMessage t;
        t <- mod_1271.get(0);
        mod_5386.put(0, t);
    endrule
    rule rule_6947;
        ChannelMessage t;
        t <- mod_3034.get(3);
        mod_5636.put(0, t);
    endrule
    rule rule_6948;
        ChannelMessage t;
        t <- mod_5309.get(121);
        mod_4961.put(0, t);
    endrule
    rule rule_6949;
        ChannelMessage t;
        t <- mod_3239.get(0);
        mod_5313.put(48, t);
    endrule
    rule rule_6950;
        ChannelMessage t;
        t <- mod_4797.get(3);
        mod_5638.put(0, t);
    endrule
    rule rule_6951;
        ChannelMessage t;
        t <- mod_1148.get(1);
        mod_5313.put(99, t);
    endrule
    rule rule_6952;
        ChannelMessage t;
        t <- mod_5394.get(0);
        mod_287.put(4, t);
    endrule
    rule rule_6953;
        ChannelMessage t;
        t <- mod_5469.get(0);
        mod_2747.put(3, t);
    endrule
    rule rule_6954;
        ChannelMessage t;
        t <- mod_4797.get(2);
        mod_5313.put(10, t);
    endrule
    rule rule_6955;
        ChannelMessage t;
        t <- mod_82.get(3);
        mod_5555.put(0, t);
    endrule
    rule rule_6956;
        ChannelMessage t;
        t <- mod_5580.get(0);
        mod_5309.put(0, t);
    endrule
    rule rule_6957;
        ChannelMessage t;
        t <- mod_2255.get(3);
        mod_5563.put(0, t);
    endrule
    rule rule_6958;
        ChannelMessage t;
        t <- mod_5254.get(0);
        mod_287.put(3, t);
    endrule
    rule rule_6959;
        ChannelMessage t;
        t <- mod_5166.get(1);
        mod_5640.put(0, t);
    endrule
    rule rule_6960;
        ChannelMessage t;
        t <- mod_5516.get(0);
        mod_2583.put(4, t);
    endrule
    rule rule_6961;
        ChannelMessage t;
        t <- mod_5600.get(34);
        mod_1394.put(1, t);
    endrule
    rule rule_6962;
        ChannelMessage t;
        t <- mod_4305.get(2);
        mod_5313.put(22, t);
    endrule
    rule rule_6963;
        ChannelMessage t;
        t <- mod_5378.get(0);
        mod_2952.put(3, t);
    endrule
    rule rule_6964;
        ChannelMessage t;
        t <- mod_5600.get(83);
        mod_3403.put(1, t);
    endrule
    rule rule_6965;
        ChannelMessage t;
        t <- mod_4756.get(2);
        mod_5313.put(11, t);
    endrule
    rule rule_6966;
        ChannelMessage t;
        t <- mod_5459.get(0);
        mod_4223.put(2, t);
    endrule
    rule rule_6967;
        ChannelMessage t;
        t <- mod_1599.get(1);
        mod_5578.put(0, t);
    endrule
    rule rule_6968;
        ChannelMessage t;
        t <- mod_779.get(2);
        mod_5484.put(0, t);
    endrule
    rule rule_6969;
        ChannelMessage t;
        t <- mod_5309.get(12);
        mod_492.put(0, t);
    endrule
    rule rule_6970;
        ChannelMessage t;
        t <- mod_738.get(1);
        mod_5307.put(0, t);
    endrule
    rule rule_6971;
        ChannelMessage t;
        t <- mod_5543.get(0);
        mod_3116.put(2, t);
    endrule
    rule rule_6972;
        ChannelMessage t;
        t <- mod_5463.get(0);
        mod_3526.put(2, t);
    endrule
    rule rule_6973;
        ChannelMessage t;
        t <- mod_4387.get(0);
        mod_5263.put(0, t);
    endrule
    rule rule_6974;
        ChannelMessage t;
        t <- mod_5600.get(74);
        mod_3034.put(1, t);
    endrule
    rule rule_6975;
        ChannelMessage t;
        t <- mod_5314.get(0);
        mod_1517.put(4, t);
    endrule
    rule rule_6976;
        ChannelMessage t;
        t <- mod_5318.get(0);
        mod_2173.put(4, t);
    endrule
    rule rule_6977;
        ChannelMessage t;
        t <- mod_4592.get(2);
        mod_5539.put(0, t);
    endrule
    rule rule_6978;
        ChannelMessage t;
        t <- mod_5302.get(0);
        mod_3362.put(4, t);
    endrule
    rule rule_6979;
        ChannelMessage t;
        t <- mod_1968.get(1);
        mod_5582.put(0, t);
    endrule
    rule rule_6980;
        ChannelMessage t;
        t <- mod_4961.get(1);
        mod_5357.put(0, t);
    endrule
    rule rule_6981;
        ChannelMessage t;
        t <- mod_5332.get(0);
        mod_1107.put(3, t);
    endrule
    rule rule_6982;
        ChannelMessage t;
        t <- mod_5338.get(0);
        mod_2460.put(4, t);
    endrule
    rule rule_6983;
        ChannelMessage t;
        t <- mod_5252.get(0);
        mod_3034.put(3, t);
    endrule
    rule rule_6984;
        ChannelMessage t;
        t <- mod_2706.get(1);
        mod_5268.put(0, t);
    endrule
    rule rule_6985;
        ChannelMessage t;
        t <- mod_5626.get(0);
        mod_5207.put(4, t);
    endrule
    rule rule_6986;
        ChannelMessage t;
        t <- mod_1230.get(1);
        mod_5465.put(0, t);
    endrule
    rule rule_6987;
        ChannelMessage t;
        t <- mod_902.get(1);
        mod_5313.put(105, t);
    endrule
    rule rule_6988;
        ChannelMessage t;
        t <- mod_492.get(1);
        mod_5477.put(0, t);
    endrule
    rule rule_6989;
        ChannelMessage t;
        t <- mod_5510.get(0);
        mod_2173.put(2, t);
    endrule
    rule rule_6990;
        ChannelMessage t;
        t <- mod_5600.get(0);
        mod_0.put(1, t);
    endrule
    rule rule_6991;
        ChannelMessage t;
        t <- mod_164.get(2);
        mod_5566.put(0, t);
    endrule
    rule rule_6992;
        ChannelMessage t;
        t <- mod_5600.get(40);
        mod_1640.put(1, t);
    endrule
    rule rule_6993;
        ChannelMessage t;
        t <- mod_1845.get(2);
        mod_5411.put(0, t);
    endrule
    rule rule_6994;
        ChannelMessage t;
        t <- mod_3116.get(1);
        mod_5470.put(0, t);
    endrule
    rule rule_6995;
        ChannelMessage t;
        t <- mod_2419.get(0);
        mod_5537.put(0, t);
    endrule
    rule rule_6996;
        ChannelMessage t;
        t <- mod_5309.get(27);
        mod_1107.put(0, t);
    endrule
    rule rule_6997;
        ChannelMessage t;
        t <- mod_3403.get(1);
        mod_5313.put(44, t);
    endrule
    rule rule_6998;
        ChannelMessage t;
        t <- mod_5370.get(0);
        mod_656.put(3, t);
    endrule
    rule rule_6999;
        ChannelMessage t;
        t <- mod_5002.get(0);
        mod_5313.put(5, t);
    endrule
    rule rule_7000;
        ChannelMessage t;
        t <- mod_5599.get(0);
        mod_369.put(4, t);
    endrule
    rule rule_7001;
        ChannelMessage t;
        t <- mod_2829.get(3);
        mod_5287.put(0, t);
    endrule
    rule rule_7002;
        ChannelMessage t;
        t <- mod_4264.get(2);
        mod_5389.put(0, t);
    endrule
    rule rule_7003;
        ChannelMessage t;
        t <- mod_4428.get(3);
        mod_5633.put(0, t);
    endrule
    rule rule_7004;
        ChannelMessage t;
        t <- mod_451.get(3);
        mod_5473.put(0, t);
    endrule
    rule rule_7005;
        ChannelMessage t;
        t <- mod_5600.get(27);
        mod_1107.put(1, t);
    endrule
    rule rule_7006;
        ChannelMessage t;
        t <- mod_5600.get(56);
        mod_2296.put(1, t);
    endrule
    rule rule_7007;
        ChannelMessage t;
        t <- mod_984.get(1);
        mod_5335.put(0, t);
    endrule
    rule rule_7008;
        ChannelMessage t;
        t <- mod_5591.get(0);
        mod_2829.put(3, t);
    endrule
    rule rule_7009;
        ChannelMessage t;
        t <- mod_5522.get(0);
        mod_2337.put(3, t);
    endrule
    rule rule_7010;
        ChannelMessage t;
        t <- mod_3526.get(1);
        mod_5463.put(0, t);
    endrule
    rule rule_7011;
        ChannelMessage t;
        t <- mod_4223.get(0);
        mod_5459.put(0, t);
    endrule
    rule rule_7012;
        ChannelMessage t;
        t <- mod_5309.get(32);
        mod_1312.put(0, t);
    endrule
    rule rule_7013;
        ChannelMessage t;
        t <- mod_5309.get(35);
        mod_1435.put(0, t);
    endrule
    rule rule_7014;
        ChannelMessage t;
        t <- mod_5371.get(0);
        mod_2296.put(2, t);
    endrule
    rule rule_7015;
        ChannelMessage t;
        t <- mod_5428.get(0);
        mod_779.put(2, t);
    endrule
    rule rule_7016;
        ChannelMessage t;
        t <- mod_5593.get(0);
        mod_3854.put(2, t);
    endrule
    rule rule_7017;
        ChannelMessage t;
        t <- mod_5278.get(0);
        mod_4756.put(2, t);
    endrule
    rule rule_7018;
        ChannelMessage t;
        t <- mod_5576.get(0);
        mod_3321.put(2, t);
    endrule
    rule rule_7019;
        ChannelMessage t;
        t <- mod_5309.get(4);
        mod_164.put(0, t);
    endrule
    rule rule_7020;
        ChannelMessage t;
        t <- mod_5600.get(108);
        mod_4428.put(1, t);
    endrule
    rule rule_7021;
        ChannelMessage t;
        t <- mod_287.get(3);
        mod_5254.put(0, t);
    endrule
    rule rule_7022;
        ChannelMessage t;
        t <- mod_2747.get(0);
        mod_5313.put(60, t);
    endrule
    rule rule_7023;
        ChannelMessage t;
        t <- mod_5528.get(0);
        mod_0.put(4, t);
    endrule
    rule rule_7024;
        ChannelMessage t;
        t <- mod_5555.get(0);
        mod_82.put(4, t);
    endrule
    rule rule_7025;
        ChannelMessage t;
        t <- mod_5396.get(0);
        mod_4797.put(3, t);
    endrule
    rule rule_7026;
        ChannelMessage t;
        t <- mod_4100.get(3);
        mod_5352.put(0, t);
    endrule
    rule rule_7027;
        ChannelMessage t;
        t <- mod_5600.get(13);
        mod_533.put(1, t);
    endrule
    rule rule_7028;
        ChannelMessage t;
        t <- mod_246.get(3);
        mod_5461.put(0, t);
    endrule
    rule rule_7029;
        ChannelMessage t;
        t <- mod_3444.get(3);
        mod_5494.put(0, t);
    endrule
    rule rule_7030;
        ChannelMessage t;
        t <- mod_2378.get(1);
        mod_5462.put(0, t);
    endrule
    rule rule_7031;
        ChannelMessage t;
        t <- mod_3854.get(2);
        mod_5322.put(0, t);
    endrule
    rule rule_7032;
        ChannelMessage t;
        t <- mod_3362.get(2);
        mod_5313.put(45, t);
    endrule
    rule rule_7033;
        ChannelMessage t;
        t <- mod_5281.get(0);
        mod_3321.put(3, t);
    endrule
    rule rule_7034;
        ChannelMessage t;
        t <- mod_492.get(2);
        mod_5404.put(0, t);
    endrule
    rule rule_7035;
        ChannelMessage t;
        t <- mod_5644.get(0);
        mod_1148.put(2, t);
    endrule
    rule rule_7036;
        ChannelMessage t;
        t <- mod_5282.get(0);
        mod_1640.put(3, t);
    endrule
    rule rule_7037;
        ChannelMessage t;
        t <- mod_3690.get(3);
        mod_5292.put(0, t);
    endrule
    rule rule_7038;
        ChannelMessage t;
        t <- mod_4469.get(0);
        mod_5300.put(0, t);
    endrule
    rule rule_7039;
        ChannelMessage t;
        t <- mod_3239.get(1);
        mod_5534.put(0, t);
    endrule
    rule rule_7040;
        ChannelMessage t;
        t <- mod_3649.get(0);
        mod_5501.put(0, t);
    endrule
    rule rule_7041;
        ChannelMessage t;
        t <- mod_5207.get(2);
        mod_5626.put(0, t);
    endrule
    rule rule_7042;
        ChannelMessage t;
        t <- mod_1599.get(2);
        mod_5257.put(0, t);
    endrule
    rule rule_7043;
        ChannelMessage t;
        t <- mod_5309.get(36);
        mod_1476.put(0, t);
    endrule
    rule rule_7044;
        ChannelMessage t;
        t <- mod_5513.get(0);
        mod_1353.put(2, t);
    endrule
    rule rule_7045;
        ChannelMessage t;
        t <- mod_5600.get(11);
        mod_451.put(1, t);
    endrule
    rule rule_7046;
        ChannelMessage t;
        t <- mod_5477.get(0);
        mod_492.put(3, t);
    endrule
    rule rule_7047;
        ChannelMessage t;
        t <- mod_5600.get(31);
        mod_1271.put(1, t);
    endrule
    rule rule_7048;
        ChannelMessage t;
        t <- mod_2173.get(2);
        mod_5318.put(0, t);
    endrule
    rule rule_7049;
        ChannelMessage t;
        t <- mod_3854.get(0);
        mod_5506.put(0, t);
    endrule
    rule rule_7050;
        ChannelMessage t;
        t <- mod_328.get(2);
        mod_5311.put(0, t);
    endrule
    rule rule_7051;
        ChannelMessage t;
        t <- mod_4182.get(3);
        mod_5609.put(0, t);
    endrule
    rule rule_7052;
        ChannelMessage t;
        t <- mod_5125.get(1);
        mod_5632.put(0, t);
    endrule
    rule rule_7053;
        ChannelMessage t;
        t <- mod_5358.get(0);
        mod_123.put(4, t);
    endrule
    rule rule_7054;
        ChannelMessage t;
        t <- mod_861.get(2);
        mod_5433.put(0, t);
    endrule
    rule rule_7055;
        ChannelMessage t;
        t <- mod_5309.get(85);
        mod_3485.put(0, t);
    endrule
    rule rule_7056;
        ChannelMessage t;
        t <- mod_5331.get(0);
        mod_1271.put(2, t);
    endrule
    rule rule_7057;
        ChannelMessage t;
        t <- mod_5393.get(0);
        mod_1312.put(4, t);
    endrule
    rule rule_7058;
        ChannelMessage t;
        t <- mod_5600.get(114);
        mod_4674.put(1, t);
    endrule
    rule rule_7059;
        ChannelMessage t;
        t <- mod_1804.get(0);
        mod_5277.put(0, t);
    endrule
    rule rule_7060;
        ChannelMessage t;
        t <- mod_1927.get(0);
        mod_5305.put(0, t);
    endrule
    rule rule_7061;
        ChannelMessage t;
        t <- mod_4592.get(1);
        mod_5427.put(0, t);
    endrule
    rule rule_7062;
        ChannelMessage t;
        t <- mod_5276.get(0);
        mod_4920.put(4, t);
    endrule
    rule rule_7063;
        ChannelMessage t;
        t <- mod_5309.get(120);
        mod_4920.put(0, t);
    endrule
    rule rule_7064;
        ChannelMessage t;
        t <- mod_5600.get(123);
        mod_5043.put(1, t);
    endrule
    rule rule_7065;
        ChannelMessage t;
        t <- mod_1476.get(2);
        mod_5581.put(0, t);
    endrule
    rule rule_7066;
        ChannelMessage t;
        t <- mod_4756.get(3);
        mod_5616.put(0, t);
    endrule
    rule rule_7067;
        ChannelMessage t;
        t <- mod_5309.get(20);
        mod_820.put(0, t);
    endrule
    rule rule_7068;
        ChannelMessage t;
        t <- mod_5309.get(98);
        mod_4018.put(0, t);
    endrule
    rule rule_7069;
        ChannelMessage t;
        t <- mod_5600.get(96);
        mod_3936.put(1, t);
    endrule
    rule rule_7070;
        ChannelMessage t;
        t <- mod_5309.get(94);
        mod_3854.put(0, t);
    endrule
    rule rule_7071;
        ChannelMessage t;
        t <- mod_5586.get(0);
        mod_3280.put(4, t);
    endrule
    rule rule_7072;
        ChannelMessage t;
        t <- mod_369.get(0);
        mod_5424.put(0, t);
    endrule
    rule rule_7073;
        ChannelMessage t;
        t <- mod_5600.get(76);
        mod_3116.put(1, t);
    endrule
    rule rule_7074;
        ChannelMessage t;
        t <- mod_5600.get(112);
        mod_4592.put(1, t);
    endrule
    rule rule_7075;
        ChannelMessage t;
        t <- mod_3280.get(1);
        mod_5295.put(0, t);
    endrule
    rule rule_7076;
        ChannelMessage t;
        t <- mod_5296.get(0);
        mod_984.put(4, t);
    endrule
    rule rule_7077;
        ChannelMessage t;
        t <- mod_2788.get(1);
        mod_5313.put(59, t);
    endrule
    rule rule_7078;
        ChannelMessage t;
        t <- mod_5600.get(82);
        mod_3362.put(1, t);
    endrule
    rule rule_7079;
        ChannelMessage t;
        t <- mod_5309.get(64);
        mod_2624.put(0, t);
    endrule
    rule rule_7080;
        ChannelMessage t;
        t <- mod_2009.get(2);
        mod_5313.put(78, t);
    endrule
    rule rule_7081;
        ChannelMessage t;
        t <- mod_3977.get(0);
        mod_5625.put(0, t);
    endrule
    rule rule_7082;
        ChannelMessage t;
        t <- mod_5512.get(0);
        mod_4387.put(2, t);
    endrule
    rule rule_7083;
        ChannelMessage t;
        t <- mod_615.get(0);
        mod_5343.put(0, t);
    endrule
    rule rule_7084;
        ChannelMessage t;
        t <- mod_5345.get(0);
        mod_3813.put(4, t);
    endrule
    rule rule_7085;
        ChannelMessage t;
        t <- mod_4961.get(2);
        mod_5313.put(6, t);
    endrule
    rule rule_7086;
        ChannelMessage t;
        t <- mod_5291.get(0);
        mod_2132.put(2, t);
    endrule
    rule rule_7087;
        ChannelMessage t;
        t <- mod_2501.get(2);
        mod_5541.put(0, t);
    endrule
    rule rule_7088;
        ChannelMessage t;
        t <- mod_2911.get(3);
        mod_5518.put(0, t);
    endrule
    rule rule_7089;
        ChannelMessage t;
        t <- mod_1640.get(2);
        mod_5527.put(0, t);
    endrule
    rule rule_7090;
        ChannelMessage t;
        t <- mod_1230.get(3);
        mod_5313.put(97, t);
    endrule
    rule rule_7091;
        ChannelMessage t;
        t <- mod_5273.get(0);
        mod_2788.put(4, t);
    endrule
    rule rule_7092;
        ChannelMessage t;
        t <- mod_5600.get(44);
        mod_1804.put(1, t);
    endrule
    rule rule_7093;
        ChannelMessage t;
        t <- mod_1886.get(2);
        mod_5313.put(81, t);
    endrule
    rule rule_7094;
        ChannelMessage t;
        t <- mod_5415.get(0);
        mod_2993.put(3, t);
    endrule
    rule rule_7095;
        ChannelMessage t;
        t <- mod_5529.get(0);
        mod_5084.put(3, t);
    endrule
    rule rule_7096;
        ChannelMessage t;
        t <- mod_3895.get(1);
        mod_5313.put(32, t);
    endrule
    rule rule_7097;
        ChannelMessage t;
        t <- mod_5334.get(0);
        mod_943.put(2, t);
    endrule
    rule rule_7098;
        ChannelMessage t;
        t <- mod_5294.get(0);
        mod_4920.put(2, t);
    endrule
    rule rule_7099;
        ChannelMessage t;
        t <- mod_3198.get(1);
        mod_5383.put(0, t);
    endrule
    rule rule_7100;
        ChannelMessage t;
        t <- mod_5320.get(0);
        mod_4674.put(4, t);
    endrule
    rule rule_7101;
        ChannelMessage t;
        t <- mod_5309.get(105);
        mod_4305.put(0, t);
    endrule
    rule rule_7102;
        ChannelMessage t;
        t <- mod_5292.get(0);
        mod_3690.put(3, t);
    endrule
    rule rule_7103;
        ChannelMessage t;
        t <- mod_1681.get(0);
        mod_5568.put(0, t);
    endrule
    rule rule_7104;
        ChannelMessage t;
        t <- mod_1107.get(2);
        mod_5434.put(0, t);
    endrule
    rule rule_7105;
        ChannelMessage t;
        t <- mod_656.get(0);
        mod_5313.put(111, t);
    endrule
    rule rule_7106;
        ChannelMessage t;
        t <- mod_3977.get(1);
        mod_5313.put(30, t);
    endrule
    rule rule_7107;
        ChannelMessage t;
        t <- mod_3444.get(1);
        mod_5313.put(43, t);
    endrule
    rule rule_7108;
        ChannelMessage t;
        t <- mod_5637.get(0);
        mod_3034.put(2, t);
    endrule
    rule rule_7109;
        ChannelMessage t;
        t <- mod_246.get(1);
        mod_5313.put(121, t);
    endrule
    rule rule_7110;
        ChannelMessage t;
        t <- mod_5600.get(125);
        mod_5125.put(1, t);
    endrule
    rule rule_7111;
        ChannelMessage t;
        t <- mod_5487.get(0);
        mod_3731.put(4, t);
    endrule
    rule rule_7112;
        ChannelMessage t;
        t <- mod_5600.get(84);
        mod_3444.put(1, t);
    endrule
    rule rule_7113;
        ChannelMessage t;
        t <- mod_5309.get(7);
        mod_287.put(0, t);
    endrule
    rule rule_7114;
        ChannelMessage t;
        t <- mod_3280.get(3);
        mod_5556.put(0, t);
    endrule
    rule rule_7115;
        ChannelMessage t;
        t <- mod_2132.get(2);
        mod_5533.put(0, t);
    endrule
    rule rule_7116;
        ChannelMessage t;
        t <- mod_205.get(3);
        mod_5359.put(0, t);
    endrule
    rule rule_7117;
        ChannelMessage t;
        t <- mod_451.get(1);
        mod_5480.put(0, t);
    endrule
    rule rule_7118;
        ChannelMessage t;
        t <- mod_3485.get(1);
        mod_5618.put(0, t);
    endrule
    rule rule_7119;
        ChannelMessage t;
        t <- mod_984.get(2);
        mod_5296.put(0, t);
    endrule
    rule rule_7120;
        ChannelMessage t;
        t <- mod_2870.get(2);
        mod_5435.put(0, t);
    endrule
    rule rule_7121;
        ChannelMessage t;
        t <- mod_5600.get(95);
        mod_3895.put(1, t);
    endrule
    rule rule_7122;
        ChannelMessage t;
        t <- mod_2624.get(2);
        mod_5615.put(0, t);
    endrule
    rule rule_7123;
        ChannelMessage t;
        t <- mod_5641.get(0);
        mod_3321.put(4, t);
    endrule
    rule rule_7124;
        ChannelMessage t;
        t <- mod_369.get(3);
        mod_5313.put(118, t);
    endrule
    rule rule_7125;
        ChannelMessage t;
        t <- mod_5309.get(10);
        mod_410.put(0, t);
    endrule
    rule rule_7126;
        ChannelMessage t;
        t <- mod_4592.get(0);
        mod_5313.put(15, t);
    endrule
    rule rule_7127;
        ChannelMessage t;
        t <- mod_4879.get(2);
        mod_5313.put(8, t);
    endrule
    rule rule_7128;
        ChannelMessage t;
        t <- mod_5043.get(1);
        mod_5486.put(0, t);
    endrule
    rule rule_7129;
        ChannelMessage t;
        t <- mod_5309.get(43);
        mod_1763.put(0, t);
    endrule
    rule rule_7130;
        ChannelMessage t;
        t <- mod_533.get(3);
        mod_5313.put(114, t);
    endrule
    rule rule_7131;
        ChannelMessage t;
        t <- mod_697.get(3);
        mod_5313.put(110, t);
    endrule
    rule rule_7132;
        ChannelMessage t;
        t <- mod_5600.get(46);
        mod_1886.put(1, t);
    endrule
    rule rule_7133;
        ChannelMessage t;
        t <- mod_5308.get(0);
        mod_1066.put(4, t);
    endrule
    rule rule_7134;
        ChannelMessage t;
        t <- mod_5601.get(0);
        mod_656.put(2, t);
    endrule
    rule rule_7135;
        ChannelMessage t;
        t <- mod_5605.get(0);
        mod_2419.put(4, t);
    endrule
    rule rule_7136;
        ChannelMessage t;
        t <- mod_4223.get(3);
        mod_5643.put(0, t);
    endrule
    rule rule_7137;
        ChannelMessage t;
        t <- mod_4961.get(3);
        mod_5505.put(0, t);
    endrule
    rule rule_7138;
        ChannelMessage t;
        t <- mod_5600.get(78);
        mod_3198.put(1, t);
    endrule
    rule rule_7139;
        ChannelMessage t;
        t <- mod_5600.get(66);
        mod_2706.put(1, t);
    endrule
    rule rule_7140;
        ChannelMessage t;
        t <- mod_5303.get(0);
        mod_3608.put(3, t);
    endrule
    rule rule_7141;
        ChannelMessage t;
        t <- mod_5600.get(92);
        mod_3772.put(1, t);
    endrule
    rule rule_7142;
        ChannelMessage t;
        t <- mod_5424.get(0);
        mod_369.put(2, t);
    endrule
    rule rule_7143;
        ChannelMessage t;
        t <- mod_5454.get(0);
        mod_2870.put(3, t);
    endrule
    rule rule_7144;
        ChannelMessage t;
        t <- mod_1435.get(1);
        mod_5367.put(0, t);
    endrule
    rule rule_7145;
        ChannelMessage t;
        t <- mod_2419.get(1);
        mod_5444.put(0, t);
    endrule
    rule rule_7146;
        ChannelMessage t;
        t <- mod_2993.get(3);
        mod_5412.put(0, t);
    endrule
    rule rule_7147;
        ChannelMessage t;
        t <- mod_3526.get(3);
        mod_5603.put(0, t);
    endrule
    rule rule_7148;
        ChannelMessage t;
        t <- mod_3567.get(3);
        mod_5315.put(0, t);
    endrule
    rule rule_7149;
        ChannelMessage t;
        t <- mod_5505.get(0);
        mod_4961.put(4, t);
    endrule
    rule rule_7150;
        ChannelMessage t;
        t <- mod_5309.get(59);
        mod_2419.put(0, t);
    endrule
    rule rule_7151;
        ChannelMessage t;
        t <- mod_3772.get(3);
        mod_5612.put(0, t);
    endrule
    rule rule_7152;
        ChannelMessage t;
        t <- mod_1968.get(0);
        mod_5313.put(79, t);
    endrule
    rule rule_7153;
        ChannelMessage t;
        t <- mod_5309.get(28);
        mod_1148.put(0, t);
    endrule
    rule rule_7154;
        ChannelMessage t;
        t <- mod_820.get(1);
        mod_5339.put(0, t);
    endrule
    rule rule_7155;
        ChannelMessage t;
        t <- mod_5600.get(6);
        mod_246.put(1, t);
    endrule
    rule rule_7156;
        ChannelMessage t;
        t <- mod_5600.get(16);
        mod_656.put(1, t);
    endrule
    rule rule_7157;
        ChannelMessage t;
        t <- mod_5600.get(39);
        mod_1599.put(1, t);
    endrule
    rule rule_7158;
        ChannelMessage t;
        t <- mod_492.get(0);
        mod_5313.put(115, t);
    endrule
    rule rule_7159;
        ChannelMessage t;
        t <- mod_5166.get(3);
        mod_5646.put(0, t);
    endrule
    rule rule_7160;
        ChannelMessage t;
        t <- mod_5316.get(0);
        mod_533.put(4, t);
    endrule
    rule rule_7161;
        ChannelMessage t;
        t <- mod_5484.get(0);
        mod_779.put(4, t);
    endrule
    rule rule_7162;
        ChannelMessage t;
        t <- mod_5309.get(80);
        mod_3280.put(0, t);
    endrule
    rule rule_7163;
        ChannelMessage t;
        t <- mod_5456.get(0);
        mod_1640.put(2, t);
    endrule
    rule rule_7164;
        ChannelMessage t;
        t <- mod_5442.get(0);
        mod_4592.put(2, t);
    endrule
    rule rule_7165;
        ChannelMessage t;
        t <- mod_3813.get(0);
        mod_5319.put(0, t);
    endrule
    rule rule_7166;
        ChannelMessage t;
        t <- mod_2255.get(0);
        mod_5379.put(0, t);
    endrule
    rule rule_7167;
        ChannelMessage t;
        t <- mod_5309.get(86);
        mod_3526.put(0, t);
    endrule
    rule rule_7168;
        ChannelMessage t;
        t <- mod_2501.get(1);
        mod_5313.put(66, t);
    endrule
    rule rule_7169;
        ChannelMessage t;
        t <- mod_5309.get(30);
        mod_1230.put(0, t);
    endrule
    rule rule_7170;
        ChannelMessage t;
        t <- mod_5439.get(0);
        mod_4346.put(4, t);
    endrule
    rule rule_7171;
        ChannelMessage t;
        t <- mod_5285.get(0);
        mod_861.put(4, t);
    endrule
    rule rule_7172;
        ChannelMessage t;
        t <- mod_410.get(0);
        mod_5267.put(0, t);
    endrule
    rule rule_7173;
        ChannelMessage t;
        t <- mod_5600.get(77);
        mod_3157.put(1, t);
    endrule
    rule rule_7174;
        ChannelMessage t;
        t <- mod_1025.get(0);
        mod_5624.put(0, t);
    endrule
    rule rule_7175;
        ChannelMessage t;
        t <- mod_5607.get(0);
        mod_3690.put(2, t);
    endrule
    rule rule_7176;
        ChannelMessage t;
        t <- mod_5309.get(57);
        mod_2337.put(0, t);
    endrule
    rule rule_7177;
        ChannelMessage t;
        t <- mod_5606.get(0);
        mod_3567.put(3, t);
    endrule
    rule rule_7178;
        ChannelMessage t;
        t <- mod_5520.get(0);
        mod_4346.put(3, t);
    endrule
    rule rule_7179;
        ChannelMessage t;
        t <- mod_3321.get(3);
        mod_5576.put(0, t);
    endrule
    rule rule_7180;
        ChannelMessage t;
        t <- mod_5638.get(0);
        mod_4797.put(2, t);
    endrule
    rule rule_7181;
        ChannelMessage t;
        t <- mod_2296.get(0);
        mod_5313.put(71, t);
    endrule
    rule rule_7182;
        ChannelMessage t;
        t <- mod_2255.get(2);
        mod_5313.put(72, t);
    endrule
    rule rule_7183;
        ChannelMessage t;
        t <- mod_5309.get(88);
        mod_3608.put(0, t);
    endrule
    rule rule_7184;
        ChannelMessage t;
        t <- mod_4059.get(1);
        mod_5313.put(28, t);
    endrule
    rule rule_7185;
        ChannelMessage t;
        t <- mod_2870.get(0);
        mod_5313.put(57, t);
    endrule
    rule rule_7186;
        ChannelMessage t;
        t <- mod_5431.get(0);
        mod_41.put(3, t);
    endrule
    rule rule_7187;
        ChannelMessage t;
        t <- mod_3403.get(2);
        mod_5504.put(0, t);
    endrule
    rule rule_7188;
        ChannelMessage t;
        t <- mod_2993.get(2);
        mod_5258.put(0, t);
    endrule
    rule rule_7189;
        ChannelMessage t;
        t <- mod_205.get(0);
        mod_5341.put(0, t);
    endrule
    rule rule_7190;
        ChannelMessage t;
        t <- mod_5309.get(47);
        mod_1927.put(0, t);
    endrule
    rule rule_7191;
        ChannelMessage t;
        t <- mod_5295.get(0);
        mod_3280.put(2, t);
    endrule
    rule rule_7192;
        ChannelMessage t;
        t <- mod_656.get(3);
        mod_5601.put(0, t);
    endrule
    rule rule_7193;
        ChannelMessage t;
        t <- mod_1066.get(1);
        mod_5554.put(0, t);
    endrule
    rule rule_7194;
        ChannelMessage t;
        t <- mod_533.get(0);
        mod_5557.put(0, t);
    endrule
    rule rule_7195;
        ChannelMessage t;
        t <- mod_5572.get(0);
        mod_943.put(3, t);
    endrule
    rule rule_7196;
        ChannelMessage t;
        t <- mod_5125.get(3);
        mod_5446.put(0, t);
    endrule
    rule rule_7197;
        ChannelMessage t;
        t <- mod_2624.get(0);
        mod_5324.put(0, t);
    endrule
    rule rule_7198;
        ChannelMessage t;
        t <- mod_5309.get(110);
        mod_4510.put(0, t);
    endrule
    rule rule_7199;
        ChannelMessage t;
        t <- mod_5377.get(0);
        mod_5600.put(1, t);
    endrule
    rule rule_7200;
        ChannelMessage t;
        t <- mod_4141.get(0);
        mod_5467.put(0, t);
    endrule
    rule rule_7201;
        ChannelMessage t;
        t <- mod_205.get(2);
        mod_5577.put(0, t);
    endrule
    rule rule_7202;
        ChannelMessage t;
        t <- mod_5309.get(56);
        mod_2296.put(0, t);
    endrule
    rule rule_7203;
        ChannelMessage t;
        t <- mod_3116.get(0);
        mod_5449.put(0, t);
    endrule
    rule rule_7204;
        ChannelMessage t;
        t <- mod_4961.get(0);
        mod_5564.put(0, t);
    endrule
    rule rule_7205;
        ChannelMessage t;
        t <- mod_5486.get(0);
        mod_5043.put(2, t);
    endrule
    rule rule_7206;
        ChannelMessage t;
        t <- mod_3649.get(1);
        mod_5491.put(0, t);
    endrule
    rule rule_7207;
        ChannelMessage t;
        t <- mod_4633.get(0);
        mod_5492.put(0, t);
    endrule
    rule rule_7208;
        ChannelMessage t;
        t <- mod_5441.get(0);
        mod_1845.put(2, t);
    endrule
    rule rule_7209;
        ChannelMessage t;
        t <- mod_5515.get(0);
        mod_2583.put(2, t);
    endrule
    rule rule_7210;
        ChannelMessage t;
        t <- mod_5615.get(0);
        mod_2624.put(3, t);
    endrule
    rule rule_7211;
        ChannelMessage t;
        t <- mod_5368.get(0);
        mod_4510.put(4, t);
    endrule
    rule rule_7212;
        ChannelMessage t;
        t <- mod_3895.get(2);
        mod_5288.put(0, t);
    endrule
    rule rule_7213;
        ChannelMessage t;
        t <- mod_1763.get(0);
        mod_5619.put(0, t);
    endrule
    rule rule_7214;
        ChannelMessage t;
        t <- mod_5521.get(0);
        mod_3649.put(2, t);
    endrule
    rule rule_7215;
        ChannelMessage t;
        t <- mod_5600.get(49);
        mod_2009.put(1, t);
    endrule
    rule rule_7216;
        ChannelMessage t;
        t <- mod_4838.get(2);
        mod_5397.put(0, t);
    endrule
    rule rule_7217;
        ChannelMessage t;
        t <- mod_5434.get(0);
        mod_1107.put(4, t);
    endrule
    rule rule_7218;
        ChannelMessage t;
        t <- mod_5489.get(0);
        mod_164.put(4, t);
    endrule
    rule rule_7219;
        ChannelMessage t;
        t <- mod_2378.get(2);
        mod_5313.put(69, t);
    endrule
    rule rule_7220;
        ChannelMessage t;
        t <- mod_5309.get(33);
        mod_1353.put(0, t);
    endrule
    rule rule_7221;
        ChannelMessage t;
        t <- mod_5372.get(0);
        mod_5326.put(0, t);
    endrule
    rule rule_7222;
        ChannelMessage t;
        t <- mod_5270.get(0);
        mod_2296.put(3, t);
    endrule
    rule rule_7223;
        ChannelMessage t;
        t <- mod_5600.get(14);
        mod_574.put(1, t);
    endrule
    rule rule_7224;
        ChannelMessage t;
        t <- mod_0.get(3);
        mod_5351.put(0, t);
    endrule
    rule rule_7225;
        ChannelMessage t;
        t <- mod_451.get(0);
        mod_5313.put(116, t);
    endrule
    rule rule_7226;
        ChannelMessage t;
        t <- mod_3362.get(0);
        mod_5323.put(0, t);
    endrule
    rule rule_7227;
        ChannelMessage t;
        t <- mod_5309.get(18);
        mod_738.put(0, t);
    endrule
    rule rule_7228;
        ChannelMessage t;
        t <- mod_5328.get(0);
        mod_123.put(2, t);
    endrule
    rule rule_7229;
        ChannelMessage t;
        t <- mod_3198.get(0);
        mod_5448.put(0, t);
    endrule
    rule rule_7230;
        ChannelMessage t;
        t <- mod_4305.get(3);
        mod_5438.put(0, t);
    endrule
    rule rule_7231;
        ChannelMessage t;
        t <- mod_2952.get(3);
        mod_5408.put(0, t);
    endrule
    rule rule_7232;
        ChannelMessage t;
        t <- mod_5309.get(5);
        mod_205.put(0, t);
    endrule
    rule rule_7233;
        ChannelMessage t;
        t <- mod_5309.get(45);
        mod_1845.put(0, t);
    endrule
    rule rule_7234;
        ChannelMessage t;
        t <- mod_5309.get(49);
        mod_2009.put(0, t);
    endrule
    rule rule_7235;
        ChannelMessage t;
        t <- mod_5595.get(0);
        mod_2665.put(4, t);
    endrule
    rule rule_7236;
        ChannelMessage t;
        t <- mod_5600.get(105);
        mod_4305.put(1, t);
    endrule
    rule rule_7237;
        ChannelMessage t;
        t <- mod_369.get(2);
        mod_5452.put(0, t);
    endrule
    rule rule_7238;
        ChannelMessage t;
        t <- mod_615.get(2);
        mod_5313.put(112, t);
    endrule
    rule rule_7239;
        ChannelMessage t;
        t <- mod_2009.get(1);
        mod_5321.put(0, t);
    endrule
    rule rule_7240;
        ChannelMessage t;
        t <- mod_5359.get(0);
        mod_205.put(3, t);
    endrule
    rule rule_7241;
        ChannelMessage t;
        t <- mod_5600.get(126);
        mod_5166.put(1, t);
    endrule
    rule rule_7242;
        ChannelMessage t;
        t <- mod_5309.get(16);
        mod_656.put(0, t);
    endrule
    rule rule_7243;
        ChannelMessage t;
        t <- mod_1271.get(3);
        mod_5313.put(96, t);
    endrule
    rule rule_7244;
        ChannelMessage t;
        t <- mod_2050.get(1);
        mod_5325.put(0, t);
    endrule
    rule rule_7245;
        ChannelMessage t;
        t <- mod_5504.get(0);
        mod_3403.put(3, t);
    endrule
    rule rule_7246;
        ChannelMessage t;
        t <- mod_123.get(2);
        mod_5358.put(0, t);
    endrule
    rule rule_7247;
        ChannelMessage t;
        t <- mod_5575.get(0);
        mod_2624.put(4, t);
    endrule
    rule rule_7248;
        ChannelMessage t;
        t <- mod_5271.get(0);
        mod_1681.put(4, t);
    endrule
    rule rule_7249;
        ChannelMessage t;
        t <- mod_2337.get(0);
        mod_5421.put(0, t);
    endrule
    rule rule_7250;
        ChannelMessage t;
        t <- mod_4551.get(3);
        mod_5313.put(16, t);
    endrule
    rule rule_7251;
        ChannelMessage t;
        t <- mod_5309.get(34);
        mod_1394.put(0, t);
    endrule
    rule rule_7252;
        ChannelMessage t;
        t <- mod_5363.get(0);
        mod_2501.put(4, t);
    endrule
    rule rule_7253;
        ChannelMessage t;
        t <- mod_5480.get(0);
        mod_451.put(3, t);
    endrule
    rule rule_7254;
        ChannelMessage t;
        t <- mod_1066.get(3);
        mod_5262.put(0, t);
    endrule
    rule rule_7255;
        ChannelMessage t;
        t <- mod_5309.get(89);
        mod_3649.put(0, t);
    endrule
    rule rule_7256;
        ChannelMessage t;
        t <- mod_5542.get(0);
        mod_1886.put(3, t);
    endrule
    rule rule_7257;
        ChannelMessage t;
        t <- mod_287.get(2);
        mod_5394.put(0, t);
    endrule
    rule rule_7258;
        ChannelMessage t;
        t <- mod_1968.get(3);
        mod_5261.put(0, t);
    endrule
    rule rule_7259;
        ChannelMessage t;
        t <- mod_5647.get(0);
        mod_3157.put(2, t);
    endrule
    rule rule_7260;
        ChannelMessage t;
        t <- mod_5600.get(9);
        mod_369.put(1, t);
    endrule
    rule rule_7261;
        ChannelMessage t;
        t <- mod_5613.get(0);
        mod_4879.put(3, t);
    endrule
    rule rule_7262;
        ChannelMessage t;
        t <- mod_2173.get(0);
        mod_5573.put(0, t);
    endrule
    rule rule_7263;
        ChannelMessage t;
        t <- mod_2173.get(1);
        mod_5510.put(0, t);
    endrule
    rule rule_7264;
        ChannelMessage t;
        t <- mod_5639.get(0);
        mod_779.put(3, t);
    endrule
    rule rule_7265;
        ChannelMessage t;
        t <- mod_5309.get(96);
        mod_3936.put(0, t);
    endrule
    rule rule_7266;
        ChannelMessage t;
        t <- mod_5556.get(0);
        mod_3280.put(3, t);
    endrule
    rule rule_7267;
        ChannelMessage t;
        t <- mod_4305.get(0);
        mod_5594.put(0, t);
    endrule
    rule rule_7268;
        ChannelMessage t;
        t <- mod_246.get(0);
        mod_5337.put(0, t);
    endrule
    rule rule_7269;
        ChannelMessage t;
        t <- mod_4469.get(3);
        mod_5275.put(0, t);
    endrule
    rule rule_7270;
        ChannelMessage t;
        t <- mod_5506.get(0);
        mod_3854.put(3, t);
    endrule
    rule rule_7271;
        ChannelMessage t;
        t <- mod_5427.get(0);
        mod_4592.put(3, t);
    endrule
    rule rule_7272;
        ChannelMessage t;
        t <- mod_5600.get(122);
        mod_5002.put(1, t);
    endrule
    rule rule_7273;
        ChannelMessage t;
        t <- mod_5309.get(26);
        mod_1066.put(0, t);
    endrule
    rule rule_7274;
        ChannelMessage t;
        t <- mod_1927.get(3);
        mod_5349.put(0, t);
    endrule
    rule rule_7275;
        ChannelMessage t;
        t <- mod_5617.get(0);
        mod_1476.put(3, t);
    endrule
    rule rule_7276;
        ChannelMessage t;
        t <- mod_2788.get(3);
        mod_5273.put(0, t);
    endrule
    rule rule_7277;
        ChannelMessage t;
        t <- mod_5309.get(119);
        mod_4879.put(0, t);
    endrule
    rule rule_7278;
        ChannelMessage t;
        t <- mod_4674.get(2);
        mod_5320.put(0, t);
    endrule
    rule rule_7279;
        ChannelMessage t;
        t <- mod_5309.get(9);
        mod_369.put(0, t);
    endrule
    rule rule_7280;
        ChannelMessage t;
        t <- mod_4264.get(1);
        mod_5437.put(0, t);
    endrule
    rule rule_7281;
        ChannelMessage t;
        t <- mod_3608.get(1);
        mod_5313.put(39, t);
    endrule
    rule rule_7282;
        ChannelMessage t;
        t <- mod_5269.get(0);
        mod_1558.put(3, t);
    endrule
    rule rule_7283;
        ChannelMessage t;
        t <- mod_5537.get(0);
        mod_2419.put(3, t);
    endrule
    rule rule_7284;
        ChannelMessage t;
        t <- mod_1394.get(0);
        mod_5313.put(93, t);
    endrule
    rule rule_7285;
        ChannelMessage t;
        t <- mod_5633.get(0);
        mod_4428.put(2, t);
    endrule
    rule rule_7286;
        ChannelMessage t;
        t <- mod_82.get(2);
        mod_5445.put(0, t);
    endrule
    rule rule_7287;
        ChannelMessage t;
        t <- mod_1353.get(3);
        mod_5313.put(94, t);
    endrule
    rule rule_7288;
        ChannelMessage t;
        t <- mod_5309.get(116);
        mod_4756.put(0, t);
    endrule
    rule rule_7289;
        ChannelMessage t;
        t <- mod_3690.get(1);
        mod_5402.put(0, t);
    endrule
    rule rule_7290;
        ChannelMessage t;
        t <- mod_5600.get(127);
        mod_5207.put(1, t);
    endrule
    rule rule_7291;
        ChannelMessage t;
        t <- mod_5388.get(0);
        mod_5002.put(2, t);
    endrule
    rule rule_7292;
        ChannelMessage t;
        t <- mod_4715.get(2);
        mod_5317.put(0, t);
    endrule
    rule rule_7293;
        ChannelMessage t;
        t <- mod_5432.get(0);
        mod_5166.put(2, t);
    endrule
    rule rule_7294;
        ChannelMessage t;
        t <- mod_1968.get(2);
        mod_5538.put(0, t);
    endrule
    rule rule_7295;
        ChannelMessage t;
        t <- mod_3772.get(2);
        mod_5430.put(0, t);
    endrule
    rule rule_7296;
        ChannelMessage t;
        t <- mod_5418.get(0);
        mod_5084.put(4, t);
    endrule
    rule rule_7297;
        ChannelMessage t;
        t <- mod_5600.get(119);
        mod_4879.put(1, t);
    endrule
    rule rule_7298;
        ChannelMessage t;
        t <- mod_1148.get(3);
        mod_5597.put(0, t);
    endrule
    rule rule_7299;
        ChannelMessage t;
        t <- mod_2829.get(1);
        mod_5313.put(58, t);
    endrule
    rule rule_7300;
        ChannelMessage t;
        t <- mod_5351.get(0);
        mod_0.put(3, t);
    endrule
    rule rule_7301;
        ChannelMessage t;
        t <- mod_5360.get(0);
        mod_246.put(4, t);
    endrule
    rule rule_7302;
        ChannelMessage t;
        t <- mod_5600.get(85);
        mod_3485.put(1, t);
    endrule
    rule rule_7303;
        ChannelMessage t;
        t <- mod_5409.get(0);
        mod_1763.put(4, t);
    endrule
    rule rule_7304;
        ChannelMessage t;
        t <- mod_5309.get(44);
        mod_1804.put(0, t);
    endrule
    rule rule_7305;
        ChannelMessage t;
        t <- mod_5449.get(0);
        mod_3116.put(3, t);
    endrule
    rule rule_7306;
        ChannelMessage t;
        t <- mod_4264.get(3);
        mod_5336.put(0, t);
    endrule
    rule rule_7307;
        ChannelMessage t;
        t <- mod_4387.get(1);
        mod_5313.put(20, t);
    endrule
    rule rule_7308;
        ChannelMessage t;
        t <- mod_3895.get(0);
        mod_5259.put(0, t);
    endrule
    rule rule_7309;
        ChannelMessage t;
        t <- mod_5600.get(2);
        mod_82.put(1, t);
    endrule
    rule rule_7310;
        ChannelMessage t;
        t <- mod_5309.get(68);
        mod_2788.put(0, t);
    endrule
    rule rule_7311;
        ChannelMessage t;
        t <- mod_1107.get(3);
        mod_5332.put(0, t);
    endrule
    rule rule_7312;
        ChannelMessage t;
        t <- mod_1640.get(3);
        mod_5282.put(0, t);
    endrule
    rule rule_7313;
        ChannelMessage t;
        t <- mod_5305.get(0);
        mod_1927.put(2, t);
    endrule
    rule rule_7314;
        ChannelMessage t;
        t <- mod_5438.get(0);
        mod_4305.put(3, t);
    endrule
    rule rule_7315;
        ChannelMessage t;
        t <- mod_5474.get(0);
        mod_615.put(3, t);
    endrule
    rule rule_7316;
        ChannelMessage t;
        t <- mod_41.get(0);
        mod_5407.put(0, t);
    endrule
    rule rule_7317;
        ChannelMessage t;
        t <- mod_2788.get(2);
        mod_5503.put(0, t);
    endrule
    rule rule_7318;
        ChannelMessage t;
        t <- mod_5395.get(0);
        mod_5207.put(2, t);
    endrule
    rule rule_7319;
        ChannelMessage t;
        t <- mod_5389.get(0);
        mod_4264.put(2, t);
    endrule
    rule rule_7320;
        ChannelMessage t;
        t <- mod_5256.get(0);
        mod_3936.put(4, t);
    endrule
    rule rule_7321;
        ChannelMessage t;
        t <- mod_5497.get(0);
        mod_2460.put(3, t);
    endrule
    rule rule_7322;
        ChannelMessage t;
        t <- mod_697.get(0);
        mod_5561.put(0, t);
    endrule
    rule rule_7323;
        ChannelMessage t;
        t <- mod_1148.get(2);
        mod_5644.put(0, t);
    endrule
    rule rule_7324;
        ChannelMessage t;
        t <- mod_5600.get(24);
        mod_984.put(1, t);
    endrule
    rule rule_7325;
        ChannelMessage t;
        t <- mod_4223.get(2);
        mod_5313.put(24, t);
    endrule
    rule rule_7326;
        ChannelMessage t;
        t <- mod_1804.get(2);
        mod_5348.put(0, t);
    endrule
    rule rule_7327;
        ChannelMessage t;
        t <- mod_4182.get(2);
        mod_5313.put(25, t);
    endrule
    rule rule_7328;
        ChannelMessage t;
        t <- mod_1640.get(1);
        mod_5456.put(0, t);
    endrule
    rule rule_7329;
        ChannelMessage t;
        t <- mod_5309.get(109);
        mod_4469.put(0, t);
    endrule
    rule rule_7330;
        ChannelMessage t;
        t <- mod_4018.get(0);
        mod_5289.put(0, t);
    endrule
    rule rule_7331;
        ChannelMessage t;
        t <- mod_5600.get(10);
        mod_410.put(1, t);
    endrule
    rule rule_7332;
        ChannelMessage t;
        t <- mod_3157.get(1);
        mod_5266.put(0, t);
    endrule
    rule rule_7333;
        ChannelMessage t;
        t <- mod_5353.get(0);
        mod_984.put(3, t);
    endrule
    rule rule_7334;
        ChannelMessage t;
        t <- mod_3321.get(2);
        mod_5281.put(0, t);
    endrule
    rule rule_7335;
        ChannelMessage t;
        t <- mod_4633.get(2);
        mod_5565.put(0, t);
    endrule
    rule rule_7336;
        ChannelMessage t;
        t <- mod_2583.get(2);
        mod_5293.put(0, t);
    endrule
    rule rule_7337;
        ChannelMessage t;
        t <- mod_1271.get(1);
        mod_5301.put(0, t);
    endrule
    rule rule_7338;
        ChannelMessage t;
        t <- mod_5290.get(0);
        mod_1763.put(3, t);
    endrule
    rule rule_7339;
        ChannelMessage t;
        t <- mod_5482.get(0);
        mod_1394.put(4, t);
    endrule
    rule rule_7340;
        ChannelMessage t;
        t <- mod_4387.get(2);
        mod_5525.put(0, t);
    endrule
    rule rule_7341;
        ChannelMessage t;
        t <- mod_5550.get(0);
        mod_451.put(2, t);
    endrule
    rule rule_7342;
        ChannelMessage t;
        t <- mod_5600.get(63);
        mod_2583.put(1, t);
    endrule
    rule rule_7343;
        ChannelMessage t;
        t <- mod_5526.get(0);
        mod_5309.put(1, t);
    endrule
    rule rule_7344;
        ChannelMessage t;
        t <- mod_5600.get(65);
        mod_2665.put(1, t);
    endrule
    rule rule_7345;
        ChannelMessage t;
        t <- mod_2911.get(2);
        mod_5333.put(0, t);
    endrule
    rule rule_7346;
        ChannelMessage t;
        t <- mod_5309.get(97);
        mod_3977.put(0, t);
    endrule
    rule rule_7347;
        ChannelMessage t;
        t <- mod_5379.get(0);
        mod_2255.put(4, t);
    endrule
    rule rule_7348;
        ChannelMessage t;
        t <- mod_5560.get(0);
        mod_4059.put(3, t);
    endrule
    rule rule_7349;
        ChannelMessage t;
        t <- mod_5600.get(53);
        mod_2173.put(1, t);
    endrule
    rule rule_7350;
        ChannelMessage t;
        t <- mod_1804.get(3);
        mod_5628.put(0, t);
    endrule
    rule rule_7351;
        ChannelMessage t;
        t <- mod_2173.get(3);
        mod_5313.put(74, t);
    endrule
    rule rule_7352;
        ChannelMessage t;
        t <- mod_1845.get(3);
        mod_5313.put(82, t);
    endrule
    rule rule_7353;
        ChannelMessage t;
        t <- mod_5485.get(0);
        mod_2747.put(4, t);
    endrule
    rule rule_7354;
        ChannelMessage t;
        t <- mod_4018.get(2);
        mod_5313.put(29, t);
    endrule
    rule rule_7355;
        ChannelMessage t;
        t <- mod_5333.get(0);
        mod_2911.put(4, t);
    endrule
    rule rule_7356;
        ChannelMessage t;
        t <- mod_5347.get(0);
        mod_656.put(4, t);
    endrule
    rule rule_7357;
        ChannelMessage t;
        t <- mod_4756.get(0);
        mod_5265.put(0, t);
    endrule
    rule rule_7358;
        ChannelMessage t;
        t <- mod_5600.get(89);
        mod_3649.put(1, t);
    endrule
    rule rule_7359;
        ChannelMessage t;
        t <- mod_5561.get(0);
        mod_697.put(3, t);
    endrule
    rule rule_7360;
        ChannelMessage t;
        t <- mod_1107.get(0);
        mod_5313.put(100, t);
    endrule
    rule rule_7361;
        ChannelMessage t;
        t <- mod_5166.get(0);
        mod_5432.put(0, t);
    endrule
    rule rule_7362;
        ChannelMessage t;
        t <- mod_2665.get(2);
        mod_5249.put(0, t);
    endrule
    rule rule_7363;
        ChannelMessage t;
        t <- mod_5544.get(0);
        mod_3895.put(4, t);
    endrule
    rule rule_7364;
        ChannelMessage t;
        t <- mod_5563.get(0);
        mod_2255.put(2, t);
    endrule
    rule rule_7365;
        ChannelMessage t;
        t <- mod_5309.get(77);
        mod_3157.put(0, t);
    endrule
    rule rule_7366;
        ChannelMessage t;
        t <- mod_5309.get(122);
        mod_5002.put(0, t);
    endrule
    rule rule_7367;
        ChannelMessage t;
        t <- mod_5381.get(0);
        mod_738.put(2, t);
    endrule
    rule rule_7368;
        ChannelMessage t;
        t <- mod_1476.get(0);
        mod_5414.put(0, t);
    endrule
    rule rule_7369;
        ChannelMessage t;
        t <- mod_5600.get(45);
        mod_1845.put(1, t);
    endrule
    rule rule_7370;
        ChannelMessage t;
        t <- mod_533.get(2);
        mod_5488.put(0, t);
    endrule
    rule rule_7371;
        ChannelMessage t;
        t <- mod_4141.get(3);
        mod_5313.put(26, t);
    endrule
    rule rule_7372;
        ChannelMessage t;
        t <- mod_3526.get(0);
        mod_5313.put(41, t);
    endrule
    rule rule_7373;
        ChannelMessage t;
        t <- mod_5293.get(0);
        mod_2583.put(3, t);
    endrule
    rule rule_7374;
        ChannelMessage t;
        t <- mod_2952.get(1);
        mod_5313.put(55, t);
    endrule
    rule rule_7375;
        ChannelMessage t;
        t <- mod_5423.get(0);
        mod_1025.put(4, t);
    endrule
    rule rule_7376;
        ChannelMessage t;
        t <- mod_5411.get(0);
        mod_1845.put(3, t);
    endrule
    rule rule_7377;
        ChannelMessage t;
        t <- mod_5382.get(0);
        mod_902.put(3, t);
    endrule
    rule rule_7378;
        ChannelMessage t;
        t <- mod_5286.get(0);
        mod_2542.put(3, t);
    endrule
    rule rule_7379;
        ChannelMessage t;
        t <- mod_5600.get(43);
        mod_1763.put(1, t);
    endrule
    rule rule_7380;
        ChannelMessage t;
        t <- mod_2296.get(2);
        mod_5551.put(0, t);
    endrule
    rule rule_7381;
        ChannelMessage t;
        t <- mod_5436.get(0);
        mod_820.put(2, t);
    endrule
    rule rule_7382;
        ChannelMessage t;
        t <- mod_1394.get(1);
        mod_5482.put(0, t);
    endrule
    rule rule_7383;
        ChannelMessage t;
        t <- mod_5361.get(0);
        mod_3813.put(3, t);
    endrule
    rule rule_7384;
        ChannelMessage t;
        t <- mod_2993.get(0);
        mod_5415.put(0, t);
    endrule
    rule rule_7385;
        ChannelMessage t;
        t <- mod_2460.get(0);
        mod_5497.put(0, t);
    endrule
    rule rule_7386;
        ChannelMessage t;
        t <- mod_246.get(2);
        mod_5360.put(0, t);
    endrule
    rule rule_7387;
        ChannelMessage t;
        t <- mod_1230.get(0);
        mod_5390.put(0, t);
    endrule
    rule rule_7388;
        ChannelMessage t;
        t <- mod_2091.get(1);
        mod_5453.put(0, t);
    endrule
    rule rule_7389;
        ChannelMessage t;
        t <- mod_4838.get(1);
        mod_5458.put(0, t);
    endrule
    rule rule_7390;
        ChannelMessage t;
        t <- mod_5313.get(0);
        mod_5372.put(0, t);
    endrule
    rule rule_7391;
        ChannelMessage t;
        t <- mod_5600.get(19);
        mod_779.put(1, t);
    endrule
    rule rule_7392;
        ChannelMessage t;
        t <- mod_5325.get(0);
        mod_2050.put(4, t);
    endrule
    rule rule_7393;
        ChannelMessage t;
        t <- mod_3444.get(2);
        mod_5508.put(0, t);
    endrule
    rule rule_7394;
        ChannelMessage t;
        t <- mod_2993.get(1);
        mod_5313.put(54, t);
    endrule
    rule rule_7395;
        ChannelMessage t;
        t <- mod_5326.get(0);
        mod_5326.put(1, t);
    endrule
    rule rule_7396;
        ChannelMessage t;
        t <- mod_5437.get(0);
        mod_4264.put(3, t);
    endrule
    rule rule_7397;
        ChannelMessage t;
        t <- mod_5530.get(0);
        mod_1230.put(2, t);
    endrule
    rule rule_7398;
        ChannelMessage t;
        t <- mod_5592.get(0);
        mod_1394.put(2, t);
    endrule
    rule rule_7399;
        ChannelMessage t;
        t <- mod_5600.get(79);
        mod_3239.put(1, t);
    endrule
    rule rule_7400;
        ChannelMessage t;
        t <- mod_5602.get(0);
        mod_1886.put(2, t);
    endrule
    rule rule_7401;
        ChannelMessage t;
        t <- mod_902.get(2);
        mod_5419.put(0, t);
    endrule
    rule rule_7402;
        ChannelMessage t;
        t <- mod_5631.get(0);
        mod_0.put(2, t);
    endrule
    rule rule_7403;
        ChannelMessage t;
        t <- mod_5249.get(0);
        mod_2665.put(2, t);
    endrule
    rule rule_7404;
        ChannelMessage t;
        t <- mod_5600.get(5);
        mod_205.put(1, t);
    endrule
    rule rule_7405;
        ChannelMessage t;
        t <- mod_738.get(3);
        mod_5313.put(109, t);
    endrule
    rule rule_7406;
        ChannelMessage t;
        t <- mod_5309.get(38);
        mod_1558.put(0, t);
    endrule
    rule rule_7407;
        ChannelMessage t;
        t <- mod_5421.get(0);
        mod_2337.put(4, t);
    endrule
    rule rule_7408;
        ChannelMessage t;
        t <- mod_2542.get(2);
        mod_5540.put(0, t);
    endrule
    rule rule_7409;
        ChannelMessage t;
        t <- mod_5348.get(0);
        mod_1804.put(2, t);
    endrule
    rule rule_7410;
        ChannelMessage t;
        t <- mod_5433.get(0);
        mod_861.put(3, t);
    endrule
    rule rule_7411;
        ChannelMessage t;
        t <- mod_4182.get(0);
        mod_5327.put(0, t);
    endrule
    rule rule_7412;
        ChannelMessage t;
        t <- mod_1271.get(2);
        mod_5331.put(0, t);
    endrule
    rule rule_7413;
        ChannelMessage t;
        t <- mod_5330.get(0);
        mod_2378.put(2, t);
    endrule
    rule rule_7414;
        ChannelMessage t;
        t <- mod_615.get(1);
        mod_5479.put(0, t);
    endrule
    rule rule_7415;
        ChannelMessage t;
        t <- mod_2091.get(3);
        mod_5403.put(0, t);
    endrule
    rule rule_7416;
        ChannelMessage t;
        t <- mod_5625.get(0);
        mod_3977.put(4, t);
    endrule
    rule rule_7417;
        ChannelMessage t;
        t <- mod_5350.get(0);
        mod_5377.put(0, t);
    endrule
    rule rule_7418;
        ChannelMessage t;
        t <- mod_820.get(0);
        mod_5436.put(0, t);
    endrule
    rule rule_7419;
        ChannelMessage t;
        t <- mod_738.get(2);
        mod_5362.put(0, t);
    endrule
    rule rule_7420;
        ChannelMessage t;
        t <- mod_1025.get(2);
        mod_5451.put(0, t);
    endrule
    rule rule_7421;
        ChannelMessage t;
        t <- mod_2378.get(0);
        mod_5365.put(0, t);
    endrule
    rule rule_7422;
        ChannelMessage t;
        t <- mod_2829.get(0);
        mod_5608.put(0, t);
    endrule
    rule rule_7423;
        ChannelMessage t;
        t <- mod_5309.get(6);
        mod_246.put(0, t);
    endrule
    rule rule_7424;
        ChannelMessage t;
        t <- mod_5251.get(0);
        mod_328.put(4, t);
    endrule
    rule rule_7425;
        ChannelMessage t;
        t <- mod_4551.get(1);
        mod_5559.put(0, t);
    endrule
    rule rule_7426;
        ChannelMessage t;
        t <- mod_779.get(1);
        mod_5428.put(0, t);
    endrule
    rule rule_7427;
        ChannelMessage t;
        t <- mod_5309.get(58);
        mod_2378.put(0, t);
    endrule
    rule rule_7428;
        ChannelMessage t;
        t <- mod_5600.get(52);
        mod_2132.put(1, t);
    endrule
    rule rule_7429;
        ChannelMessage t;
        t <- mod_5611.get(0);
        mod_1722.put(4, t);
    endrule
    rule rule_7430;
        ChannelMessage t;
        t <- mod_3567.get(1);
        mod_5313.put(40, t);
    endrule
    rule rule_7431;
        ChannelMessage t;
        t <- mod_0.get(1);
        mod_5631.put(0, t);
    endrule
    rule rule_7432;
        ChannelMessage t;
        t <- mod_2583.get(3);
        mod_5515.put(0, t);
    endrule
    rule rule_7433;
        ChannelMessage t;
        t <- mod_5268.get(0);
        mod_2706.put(3, t);
    endrule
    rule rule_7434;
        ChannelMessage t;
        t <- mod_5265.get(0);
        mod_4756.put(3, t);
    endrule
    rule rule_7435;
        ChannelMessage t;
        t <- mod_2419.get(3);
        mod_5313.put(68, t);
    endrule
    rule rule_7436;
        ChannelMessage t;
        t <- mod_2583.get(1);
        mod_5516.put(0, t);
    endrule
    rule rule_7437;
        ChannelMessage t;
        t <- mod_5258.get(0);
        mod_2993.put(4, t);
    endrule
    rule rule_7438;
        ChannelMessage t;
        t <- mod_3403.get(3);
        mod_5596.put(0, t);
    endrule
    rule rule_7439;
        ChannelMessage t;
        t <- mod_5300.get(0);
        mod_4469.put(3, t);
    endrule
    rule rule_7440;
        ChannelMessage t;
        t <- mod_2050.get(2);
        mod_5313.put(77, t);
    endrule
    rule rule_7441;
        ChannelMessage t;
        t <- mod_5539.get(0);
        mod_4592.put(4, t);
    endrule
    rule rule_7442;
        ChannelMessage t;
        t <- mod_2665.get(3);
        mod_5374.put(0, t);
    endrule
    rule rule_7443;
        ChannelMessage t;
        t <- mod_3485.get(2);
        mod_5313.put(42, t);
    endrule
    rule rule_7444;
        ChannelMessage t;
        t <- mod_5466.get(0);
        mod_3075.put(4, t);
    endrule
    rule rule_7445;
        ChannelMessage t;
        t <- mod_5519.get(0);
        mod_4018.put(3, t);
    endrule
    rule rule_7446;
        ChannelMessage t;
        t <- mod_5535.get(0);
        mod_1517.put(2, t);
    endrule
    rule rule_7447;
        ChannelMessage t;
        t <- mod_5407.get(0);
        mod_41.put(2, t);
    endrule
    rule rule_7448;
        ChannelMessage t;
        t <- mod_5450.get(0);
        mod_1722.put(3, t);
    endrule
    rule rule_7449;
        ChannelMessage t;
        t <- mod_5386.get(0);
        mod_1271.put(3, t);
    endrule
    rule rule_7450;
        ChannelMessage t;
        t <- mod_5629.get(0);
        mod_2870.put(2, t);
    endrule
    rule rule_7451;
        ChannelMessage t;
        t <- mod_205.get(1);
        mod_5313.put(122, t);
    endrule
    rule rule_7452;
        ChannelMessage t;
        t <- mod_2337.get(3);
        mod_5502.put(0, t);
    endrule
    rule rule_7453;
        ChannelMessage t;
        t <- mod_4920.get(0);
        mod_5313.put(7, t);
    endrule
    rule rule_7454;
        ChannelMessage t;
        t <- mod_5309.get(71);
        mod_2911.put(0, t);
    endrule
    rule rule_7455;
        ChannelMessage t;
        t <- mod_5493.get(0);
        mod_3977.put(2, t);
    endrule
    rule rule_7456;
        ChannelMessage t;
        t <- mod_82.get(0);
        mod_5313.put(125, t);
    endrule
    rule rule_7457;
        ChannelMessage t;
        t <- mod_5261.get(0);
        mod_1968.put(2, t);
    endrule
    rule rule_7458;
        ChannelMessage t;
        t <- mod_5299.get(0);
        mod_1107.put(2, t);
    endrule
    rule rule_7459;
        ChannelMessage t;
        t <- mod_5309.get(51);
        mod_2091.put(0, t);
    endrule
    rule rule_7460;
        ChannelMessage t;
        t <- mod_5508.get(0);
        mod_3444.put(2, t);
    endrule
    rule rule_7461;
        ChannelMessage t;
        t <- mod_4551.get(2);
        mod_5391.put(0, t);
    endrule
    rule rule_7462;
        ChannelMessage t;
        t <- mod_3977.get(2);
        mod_5478.put(0, t);
    endrule
    rule rule_7463;
        ChannelMessage t;
        t <- mod_5574.get(0);
        mod_4059.put(4, t);
    endrule
    rule rule_7464;
        ChannelMessage t;
        t <- mod_5084.get(3);
        mod_5529.put(0, t);
    endrule
    rule rule_7465;
        ChannelMessage t;
        t <- mod_2542.get(3);
        mod_5313.put(65, t);
    endrule
    rule rule_7466;
        ChannelMessage t;
        t <- mod_4018.get(3);
        mod_5519.put(0, t);
    endrule
    rule rule_7467;
        ChannelMessage t;
        t <- mod_328.get(0);
        mod_5548.put(0, t);
    endrule
    rule rule_7468;
        ChannelMessage t;
        t <- mod_4059.get(0);
        mod_5574.put(0, t);
    endrule
    rule rule_7469;
        ChannelMessage t;
        t <- mod_5309.get(92);
        mod_3772.put(0, t);
    endrule
    rule rule_7470;
        ChannelMessage t;
        t <- mod_5324.get(0);
        mod_2624.put(2, t);
    endrule
    rule rule_7471;
        ChannelMessage t;
        t <- mod_5499.get(0);
        mod_4100.put(3, t);
    endrule
    rule rule_7472;
        ChannelMessage t;
        t <- mod_1845.get(0);
        mod_5329.put(0, t);
    endrule
    rule rule_7473;
        ChannelMessage t;
        t <- mod_2132.get(0);
        mod_5571.put(0, t);
    endrule
    rule rule_7474;
        ChannelMessage t;
        t <- mod_5207.get(1);
        mod_5395.put(0, t);
    endrule
    rule rule_7475;
        ChannelMessage t;
        t <- mod_5309.get(17);
        mod_697.put(0, t);
    endrule
    rule rule_7476;
        ChannelMessage t;
        t <- mod_5339.get(0);
        mod_820.put(4, t);
    endrule
    rule rule_7477;
        ChannelMessage t;
        t <- mod_2952.get(2);
        mod_5514.put(0, t);
    endrule
    rule rule_7478;
        ChannelMessage t;
        t <- mod_5349.get(0);
        mod_1927.put(3, t);
    endrule
    rule rule_7479;
        ChannelMessage t;
        t <- mod_5533.get(0);
        mod_2132.put(3, t);
    endrule
    rule rule_7480;
        ChannelMessage t;
        t <- mod_4141.get(2);
        mod_5425.put(0, t);
    endrule
    rule rule_7481;
        ChannelMessage t;
        t <- mod_4879.get(1);
        mod_5622.put(0, t);
    endrule
    rule rule_7482;
        ChannelMessage t;
        t <- mod_5582.get(0);
        mod_1968.put(4, t);
    endrule
    rule rule_7483;
        ChannelMessage t;
        t <- mod_4305.get(1);
        mod_5413.put(0, t);
    endrule
    rule rule_7484;
        ChannelMessage t;
        t <- mod_5084.get(0);
        mod_5614.put(0, t);
    endrule
    rule rule_7485;
        ChannelMessage t;
        t <- mod_5568.get(0);
        mod_1681.put(2, t);
    endrule
    rule rule_7486;
        ChannelMessage t;
        t <- mod_5503.get(0);
        mod_2788.put(3, t);
    endrule
    rule rule_7487;
        ChannelMessage t;
        t <- mod_1681.get(1);
        mod_5271.put(0, t);
    endrule
    rule rule_7488;
        ChannelMessage t;
        t <- mod_5253.get(0);
        mod_5043.put(3, t);
    endrule
    rule rule_7489;
        ChannelMessage t;
        t <- mod_4223.get(1);
        mod_5511.put(0, t);
    endrule
    rule rule_7490;
        ChannelMessage t;
        t <- mod_5373.get(0);
        mod_4715.put(2, t);
    endrule
    rule rule_7491;
        ChannelMessage t;
        t <- mod_5404.get(0);
        mod_492.put(2, t);
    endrule
    rule rule_7492;
        ChannelMessage t;
        t <- mod_3936.get(2);
        mod_5313.put(31, t);
    endrule
    rule rule_7493;
        ChannelMessage t;
        t <- mod_5600.get(25);
        mod_1025.put(1, t);
    endrule
    rule rule_7494;
        ChannelMessage t;
        t <- mod_1312.get(1);
        mod_5304.put(0, t);
    endrule
    rule rule_7495;
        ChannelMessage t;
        t <- mod_164.get(1);
        mod_5313.put(123, t);
    endrule
    rule rule_7496;
        ChannelMessage t;
        t <- mod_2583.get(0);
        mod_5313.put(64, t);
    endrule
    rule rule_7497;
        ChannelMessage t;
        t <- mod_3034.get(2);
        mod_5637.put(0, t);
    endrule
    rule rule_7498;
        ChannelMessage t;
        t <- mod_5309.get(83);
        mod_3403.put(0, t);
    endrule
    rule rule_7499;
        ChannelMessage t;
        t <- mod_5435.get(0);
        mod_2870.put(4, t);
    endrule
    rule rule_7500;
        ChannelMessage t;
        t <- mod_3690.get(2);
        mod_5313.put(37, t);
    endrule
    rule rule_7501;
        ChannelMessage t;
        t <- mod_5376.get(0);
        mod_4469.put(2, t);
    endrule
    rule rule_7502;
        ChannelMessage t;
        t <- mod_5309.get(40);
        mod_1640.put(0, t);
    endrule
    rule rule_7503;
        ChannelMessage t;
        t <- mod_5494.get(0);
        mod_3444.put(3, t);
    endrule
    rule rule_7504;
        ChannelMessage t;
        t <- mod_5567.get(0);
        mod_4715.put(4, t);
    endrule
    rule rule_7505;
        ChannelMessage t;
        t <- mod_5600.get(61);
        mod_2501.put(1, t);
    endrule
    rule rule_7506;
        ChannelMessage t;
        t <- mod_4674.get(1);
        mod_5313.put(13, t);
    endrule
    rule rule_7507;
        ChannelMessage t;
        t <- mod_2460.get(3);
        mod_5648.put(0, t);
    endrule
    rule rule_7508;
        ChannelMessage t;
        t <- mod_1517.get(2);
        mod_5584.put(0, t);
    endrule
    rule rule_7509;
        ChannelMessage t;
        t <- mod_5600.get(12);
        mod_492.put(1, t);
    endrule
    rule rule_7510;
        ChannelMessage t;
        t <- mod_2706.get(0);
        mod_5313.put(61, t);
    endrule
    rule rule_7511;
        ChannelMessage t;
        t <- mod_5569.get(0);
        mod_2091.put(3, t);
    endrule
    rule rule_7512;
        ChannelMessage t;
        t <- mod_5309.get(42);
        mod_1722.put(0, t);
    endrule
    rule rule_7513;
        ChannelMessage t;
        t <- mod_5416.get(0);
        mod_2214.put(3, t);
    endrule
    rule rule_7514;
        ChannelMessage t;
        t <- mod_5614.get(0);
        mod_5084.put(2, t);
    endrule
    rule rule_7515;
        ChannelMessage t;
        t <- mod_5642.get(0);
        mod_3731.put(2, t);
    endrule
    rule rule_7516;
        ChannelMessage t;
        t <- mod_5344.get(0);
        mod_5248.put(0, t);
    endrule
    rule rule_7517;
        ChannelMessage t;
        t <- mod_5507.get(0);
        mod_3198.put(3, t);
    endrule
    rule rule_7518;
        ChannelMessage t;
        t <- mod_492.get(3);
        mod_5610.put(0, t);
    endrule
    rule rule_7519;
        ChannelMessage t;
        t <- mod_5002.get(3);
        mod_5552.put(0, t);
    endrule
    rule rule_7520;
        ChannelMessage t;
        t <- mod_5250.get(0);
        mod_4428.put(4, t);
    endrule
    rule rule_7521;
        ChannelMessage t;
        t <- mod_943.get(0);
        mod_5334.put(0, t);
    endrule
    rule rule_7522;
        ChannelMessage t;
        t <- mod_1558.get(1);
        mod_5313.put(89, t);
    endrule
    rule rule_7523;
        ChannelMessage t;
        t <- mod_1845.get(1);
        mod_5441.put(0, t);
    endrule
    rule rule_7524;
        ChannelMessage t;
        t <- mod_5600.get(106);
        mod_4346.put(1, t);
    endrule
    rule rule_7525;
        ChannelMessage t;
        t <- mod_5275.get(0);
        mod_4469.put(4, t);
    endrule
    rule rule_7526;
        ChannelMessage t;
        t <- mod_5632.get(0);
        mod_5125.put(3, t);
    endrule
    rule rule_7527;
        ChannelMessage t;
        t <- mod_5309.get(79);
        mod_3239.put(0, t);
    endrule
    rule rule_7528;
        ChannelMessage t;
        t <- mod_2747.get(2);
        mod_5469.put(0, t);
    endrule
    rule rule_7529;
        ChannelMessage t;
        t <- mod_4715.get(1);
        mod_5313.put(12, t);
    endrule
    rule rule_7530;
        ChannelMessage t;
        t <- mod_5366.get(0);
        mod_4059.put(2, t);
    endrule
    rule rule_7531;
        ChannelMessage t;
        t <- mod_5634.get(0);
        mod_4674.put(3, t);
    endrule
    rule rule_7532;
        ChannelMessage t;
        t <- mod_943.get(1);
        mod_5572.put(0, t);
    endrule
    rule rule_7533;
        ChannelMessage t;
        t <- mod_5623.get(0);
        mod_2050.put(3, t);
    endrule
    rule rule_7534;
        ChannelMessage t;
        t <- mod_2747.get(1);
        mod_5422.put(0, t);
    endrule
    rule rule_7535;
        ChannelMessage t;
        t <- mod_5585.get(0);
        mod_3075.put(3, t);
    endrule
    rule rule_7536;
        ChannelMessage t;
        t <- mod_5467.get(0);
        mod_4141.put(3, t);
    endrule
    rule rule_7537;
        ChannelMessage t;
        t <- mod_5554.get(0);
        mod_1066.put(3, t);
    endrule
    rule rule_7538;
        ChannelMessage t;
        t <- mod_5600.get(7);
        mod_287.put(1, t);
    endrule
    rule rule_7539;
        ChannelMessage t;
        t <- mod_410.get(2);
        mod_5604.put(0, t);
    endrule
    rule rule_7540;
        ChannelMessage t;
        t <- mod_5430.get(0);
        mod_3772.put(3, t);
    endrule
    rule rule_7541;
        ChannelMessage t;
        t <- mod_4264.get(0);
        mod_5313.put(23, t);
    endrule
    rule rule_7542;
        ChannelMessage t;
        t <- mod_5577.get(0);
        mod_205.put(2, t);
    endrule
    rule rule_7543;
        ChannelMessage t;
        t <- mod_369.get(1);
        mod_5599.put(0, t);
    endrule
    rule rule_7544;
        ChannelMessage t;
        t <- mod_1312.get(2);
        mod_5393.put(0, t);
    endrule
    rule rule_7545;
        ChannelMessage t;
        t <- mod_5600.get(30);
        mod_1230.put(1, t);
    endrule
    rule rule_7546;
        ChannelMessage t;
        t <- mod_5309.get(2);
        mod_82.put(0, t);
    endrule
    rule rule_7547;
        ChannelMessage t;
        t <- mod_5309.get(23);
        mod_943.put(0, t);
    endrule
    rule rule_7548;
        ChannelMessage t;
        t <- mod_5488.get(0);
        mod_533.put(3, t);
    endrule
    rule rule_7549;
        ChannelMessage t;
        t <- mod_451.get(2);
        mod_5550.put(0, t);
    endrule
    rule rule_7550;
        ChannelMessage t;
        t <- mod_5279.get(0);
        mod_3772.put(4, t);
    endrule
    rule rule_7551;
        ChannelMessage t;
        t <- mod_5517.get(0);
        mod_574.put(2, t);
    endrule
    rule rule_7552;
        ChannelMessage t;
        t <- mod_5479.get(0);
        mod_615.put(2, t);
    endrule
    rule rule_7553;
        ChannelMessage t;
        t <- mod_3731.get(3);
        mod_5313.put(36, t);
    endrule
    rule rule_7554;
        ChannelMessage t;
        t <- mod_5367.get(0);
        mod_1435.put(4, t);
    endrule
    rule rule_7555;
        ChannelMessage t;
        t <- mod_5600.get(113);
        mod_4633.put(1, t);
    endrule
    rule rule_7556;
        ChannelMessage t;
        t <- mod_3403.get(0);
        mod_5553.put(0, t);
    endrule
    rule rule_7557;
        ChannelMessage t;
        t <- mod_5541.get(0);
        mod_2501.put(3, t);
    endrule
    rule rule_7558;
        ChannelMessage t;
        t <- mod_2214.get(1);
        mod_5313.put(73, t);
    endrule
    rule rule_7559;
        ChannelMessage t;
        t <- mod_4797.get(1);
        mod_5396.put(0, t);
    endrule
    rule rule_7560;
        ChannelMessage t;
        t <- mod_2050.get(0);
        mod_5623.put(0, t);
    endrule
    rule rule_7561;
        ChannelMessage t;
        t <- mod_656.get(1);
        mod_5347.put(0, t);
    endrule
    rule rule_7562;
        ChannelMessage t;
        t <- mod_1558.get(3);
        mod_5589.put(0, t);
    endrule
    rule rule_7563;
        ChannelMessage t;
        t <- mod_5392.get(0);
        mod_287.put(2, t);
    endrule
    rule rule_7564;
        ChannelMessage t;
        t <- mod_5476.get(0);
        mod_3936.put(2, t);
    endrule
    rule rule_7565;
        ChannelMessage t;
        t <- mod_5612.get(0);
        mod_3772.put(2, t);
    endrule
    rule rule_7566;
        ChannelMessage t;
        t <- mod_2091.get(0);
        mod_5569.put(0, t);
    endrule
    rule rule_7567;
        ChannelMessage t;
        t <- mod_5600.get(38);
        mod_1558.put(1, t);
    endrule
    rule rule_7568;
        ChannelMessage t;
        t <- mod_1148.get(0);
        mod_5260.put(0, t);
    endrule
    rule rule_7569;
        ChannelMessage t;
        t <- mod_1517.get(1);
        mod_5314.put(0, t);
    endrule
    rule rule_7570;
        ChannelMessage t;
        t <- mod_5483.get(0);
        mod_697.put(4, t);
    endrule
    rule rule_7571;
        ChannelMessage t;
        t <- mod_5262.get(0);
        mod_1066.put(2, t);
    endrule
    rule rule_7572;
        ChannelMessage t;
        t <- mod_1189.get(0);
        mod_5387.put(0, t);
    endrule
    rule rule_7573;
        ChannelMessage t;
        t <- mod_2255.get(1);
        mod_5364.put(0, t);
    endrule
    rule rule_7574;
        ChannelMessage t;
        t <- mod_5309.get(67);
        mod_2747.put(0, t);
    endrule
    rule rule_7575;
        ChannelMessage t;
        t <- mod_287.get(1);
        mod_5392.put(0, t);
    endrule
    rule rule_7576;
        ChannelMessage t;
        t <- mod_5600.get(23);
        mod_943.put(1, t);
    endrule
    rule rule_7577;
        ChannelMessage t;
        t <- mod_3649.get(3);
        mod_5521.put(0, t);
    endrule
    rule rule_7578;
        ChannelMessage t;
        t <- mod_4920.get(1);
        mod_5276.put(0, t);
    endrule
    rule rule_7579;
        ChannelMessage t;
        t <- mod_5309.get(65);
        mod_2665.put(0, t);
    endrule
    rule rule_7580;
        ChannelMessage t;
        t <- mod_5309.get(84);
        mod_3444.put(0, t);
    endrule
    rule rule_7581;
        ChannelMessage t;
        t <- mod_5472.get(0);
        mod_164.put(2, t);
    endrule
    rule rule_7582;
        ChannelMessage t;
        t <- mod_5309.get(19);
        mod_779.put(0, t);
    endrule
    rule rule_7583;
        ChannelMessage t;
        t <- mod_5346.get(0);
        mod_3608.put(2, t);
    endrule
    rule rule_7584;
        ChannelMessage t;
        t <- mod_5417.get(0);
        mod_1435.put(2, t);
    endrule
    rule rule_7585;
        ChannelMessage t;
        t <- mod_5536.get(0);
        mod_4920.put(3, t);
    endrule
    rule rule_7586;
        ChannelMessage t;
        t <- mod_1189.get(1);
        mod_5313.put(98, t);
    endrule
    rule rule_7587;
        ChannelMessage t;
        t <- mod_5272.get(0);
        mod_82.put(3, t);
    endrule
    rule rule_7588;
        ChannelMessage t;
        t <- mod_2296.get(1);
        mod_5371.put(0, t);
    endrule
    rule rule_7589;
        ChannelMessage t;
        t <- mod_5309.get(114);
        mod_4674.put(0, t);
    endrule
    rule rule_7590;
        ChannelMessage t;
        t <- mod_1353.get(2);
        mod_5513.put(0, t);
    endrule
    rule rule_7591;
        ChannelMessage t;
        t <- mod_1722.get(2);
        mod_5313.put(85, t);
    endrule
    rule rule_7592;
        ChannelMessage t;
        t <- mod_5356.get(0);
        mod_2009.put(2, t);
    endrule
    rule rule_7593;
        ChannelMessage t;
        t <- mod_5043.get(2);
        mod_5253.put(0, t);
    endrule
    rule rule_7594;
        ChannelMessage t;
        t <- mod_5453.get(0);
        mod_2091.put(4, t);
    endrule
    rule rule_7595;
        ChannelMessage t;
        t <- mod_3034.get(0);
        mod_5313.put(53, t);
    endrule
    rule rule_7596;
        ChannelMessage t;
        t <- mod_5309.get(0);
        mod_0.put(0, t);
    endrule
    rule rule_7597;
        ChannelMessage t;
        t <- mod_5495.get(0);
        mod_5255.put(0, t);
    endrule
    rule rule_7598;
        ChannelMessage t;
        t <- mod_5559.get(0);
        mod_4551.put(4, t);
    endrule
    rule rule_7599;
        ChannelMessage t;
        t <- mod_3280.get(2);
        mod_5586.put(0, t);
    endrule
    rule rule_7600;
        ChannelMessage t;
        t <- mod_5443.get(0);
        mod_1189.put(2, t);
    endrule
    rule rule_7601;
        ChannelMessage t;
        t <- mod_5362.get(0);
        mod_738.put(3, t);
    endrule
    rule rule_7602;
        ChannelMessage t;
        t <- mod_5400.get(0);
        mod_3485.put(3, t);
    endrule
    rule rule_7603;
        ChannelMessage t;
        t <- mod_1394.get(2);
        mod_5579.put(0, t);
    endrule
    rule rule_7604;
        ChannelMessage t;
        t <- mod_5248.get(0);
        mod_5580.put(0, t);
    endrule
    rule rule_7605;
        ChannelMessage t;
        t <- mod_5259.get(0);
        mod_3895.put(2, t);
    endrule
    rule rule_7606;
        ChannelMessage t;
        t <- mod_5369.get(0);
        mod_2501.put(2, t);
    endrule
    rule rule_7607;
        ChannelMessage t;
        t <- mod_5600.get(70);
        mod_2870.put(1, t);
    endrule
    rule rule_7608;
        ChannelMessage t;
        t <- mod_5319.get(0);
        mod_3813.put(2, t);
    endrule
    rule rule_7609;
        ChannelMessage t;
        t <- mod_5600.get(111);
        mod_4551.put(1, t);
    endrule
    rule rule_7610;
        ChannelMessage t;
        t <- mod_0.get(2);
        mod_5528.put(0, t);
    endrule
    rule rule_7611;
        ChannelMessage t;
        t <- mod_5478.get(0);
        mod_3977.put(3, t);
    endrule
    rule rule_7612;
        ChannelMessage t;
        t <- mod_5616.get(0);
        mod_4756.put(4, t);
    endrule
    rule rule_7613;
        ChannelMessage t;
        t <- mod_5557.get(0);
        mod_533.put(2, t);
    endrule
    rule rule_7614;
        ChannelMessage t;
        t <- mod_5600.get(42);
        mod_1722.put(1, t);
    endrule
    rule rule_7615;
        ChannelMessage t;
        t <- mod_2214.get(0);
        mod_5416.put(0, t);
    endrule
    rule rule_7616;
        ChannelMessage t;
        t <- mod_5309.get(111);
        mod_4551.put(0, t);
    endrule
    rule rule_7617;
        ChannelMessage t;
        t <- mod_3116.get(2);
        mod_5313.put(51, t);
    endrule
    rule rule_7618;
        ChannelMessage t;
        t <- mod_3198.get(2);
        mod_5313.put(49, t);
    endrule
    rule rule_7619;
        ChannelMessage t;
        t <- mod_123.get(3);
        mod_5500.put(0, t);
    endrule
    rule rule_7620;
        ChannelMessage t;
        t <- mod_41.get(1);
        mod_5431.put(0, t);
    endrule
    rule rule_7621;
        ChannelMessage t;
        t <- mod_5548.get(0);
        mod_328.put(3, t);
    endrule
    rule rule_7622;
        ChannelMessage t;
        t <- mod_5309.get(90);
        mod_3690.put(0, t);
    endrule
    rule rule_7623;
        ChannelMessage t;
        t <- mod_287.get(0);
        mod_5313.put(120, t);
    endrule
    rule rule_7624;
        ChannelMessage t;
        t <- mod_5600.get(62);
        mod_2542.put(1, t);
    endrule
    rule rule_7625;
        ChannelMessage t;
        t <- mod_3649.get(2);
        mod_5313.put(38, t);
    endrule
    rule rule_7626;
        ChannelMessage t;
        t <- mod_656.get(2);
        mod_5370.put(0, t);
    endrule
    rule rule_7627;
        ChannelMessage t;
        t <- mod_4469.get(1);
        mod_5376.put(0, t);
    endrule
    rule rule_7628;
        ChannelMessage t;
        t <- mod_2378.get(3);
        mod_5330.put(0, t);
    endrule
    rule rule_7629;
        ChannelMessage t;
        t <- mod_5600.get(54);
        mod_2214.put(1, t);
    endrule
    rule rule_7630;
        ChannelMessage t;
        t <- mod_5354.get(0);
        mod_4797.put(4, t);
    endrule
    rule rule_7631;
        ChannelMessage t;
        t <- mod_5335.get(0);
        mod_984.put(2, t);
    endrule
    rule rule_7632;
        ChannelMessage t;
        t <- mod_5315.get(0);
        mod_3567.put(4, t);
    endrule
    rule rule_7633;
        ChannelMessage t;
        t <- mod_5309.get(53);
        mod_2173.put(0, t);
    endrule
    rule rule_7634;
        ChannelMessage t;
        t <- mod_3854.get(3);
        mod_5313.put(33, t);
    endrule
    rule rule_7635;
        ChannelMessage t;
        t <- mod_5600.get(51);
        mod_2091.put(1, t);
    endrule
    rule rule_7636;
        ChannelMessage t;
        t <- mod_5603.get(0);
        mod_3526.put(4, t);
    endrule
    rule rule_7637;
        ChannelMessage t;
        t <- mod_5452.get(0);
        mod_369.put(3, t);
    endrule
    rule rule_7638;
        ChannelMessage t;
        t <- mod_5309.get(104);
        mod_4264.put(0, t);
    endrule
    rule rule_7639;
        ChannelMessage t;
        t <- mod_5297.get(0);
        mod_2706.put(2, t);
    endrule
    rule rule_7640;
        ChannelMessage t;
        t <- mod_5600.get(58);
        mod_2378.put(1, t);
    endrule
    rule rule_7641;
        ChannelMessage t;
        t <- mod_4879.get(3);
        mod_5524.put(0, t);
    endrule
    rule rule_7642;
        ChannelMessage t;
        t <- mod_5600.get(41);
        mod_1681.put(1, t);
    endrule
    rule rule_7643;
        ChannelMessage t;
        t <- mod_1435.get(2);
        mod_5283.put(0, t);
    endrule
    rule rule_7644;
        ChannelMessage t;
        t <- mod_5309.get(14);
        mod_574.put(0, t);
    endrule
    rule rule_7645;
        ChannelMessage t;
        t <- mod_1189.get(2);
        mod_5583.put(0, t);
    endrule
    rule rule_7646;
        ChannelMessage t;
        t <- mod_5645.get(0);
        mod_2788.put(2, t);
    endrule
    rule rule_7647;
        ChannelMessage t;
        t <- mod_5309.get(61);
        mod_2501.put(0, t);
    endrule
    rule rule_7648;
        ChannelMessage t;
        t <- mod_5630.get(0);
        mod_1599.put(3, t);
    endrule
    rule rule_7649;
        ChannelMessage t;
        t <- mod_5628.get(0);
        mod_1804.put(4, t);
    endrule
    rule rule_7650;
        ChannelMessage t;
        t <- mod_2214.get(2);
        mod_5590.put(0, t);
    endrule
    rule rule_7651;
        ChannelMessage t;
        t <- mod_5534.get(0);
        mod_3239.put(2, t);
    endrule
    rule rule_7652;
        ChannelMessage t;
        t <- mod_1763.get(1);
        mod_5313.put(84, t);
    endrule
    rule rule_7653;
        ChannelMessage t;
        t <- mod_0.get(0);
        mod_5313.put(127, t);
    endrule
    rule rule_7654;
        ChannelMessage t;
        t <- mod_5600.get(98);
        mod_4018.put(1, t);
    endrule
    rule rule_7655;
        ChannelMessage t;
        t <- mod_5309.get(69);
        mod_2829.put(0, t);
    endrule
    rule rule_7656;
        ChannelMessage t;
        t <- mod_5309.get(95);
        mod_3895.put(0, t);
    endrule
    rule rule_7657;
        ChannelMessage t;
        t <- mod_2665.get(1);
        mod_5313.put(62, t);
    endrule
    rule rule_7658;
        ChannelMessage t;
        t <- mod_5471.get(0);
        mod_1353.put(4, t);
    endrule
    rule rule_7659;
        ChannelMessage t;
        t <- mod_5309.get(127);
        mod_5207.put(0, t);
    endrule
    rule rule_7660;
        ChannelMessage t;
        t <- mod_4387.get(3);
        mod_5512.put(0, t);
    endrule
    rule rule_7661;
        ChannelMessage t;
        t <- mod_2706.get(3);
        mod_5406.put(0, t);
    endrule
    rule rule_7662;
        ChannelMessage t;
        t <- mod_4510.get(2);
        mod_5509.put(0, t);
    endrule
    rule rule_7663;
        ChannelMessage t;
        t <- mod_5600.get(120);
        mod_4920.put(1, t);
    endrule
    rule rule_7664;
        ChannelMessage t;
        t <- mod_5547.get(0);
        mod_902.put(4, t);
    endrule
    rule rule_7665;
        ChannelMessage t;
        t <- mod_1640.get(0);
        mod_5313.put(87, t);
    endrule
    rule rule_7666;
        ChannelMessage t;
        t <- mod_5540.get(0);
        mod_2542.put(4, t);
    endrule
    rule rule_7667;
        ChannelMessage t;
        t <- mod_5558.get(0);
        mod_4510.put(3, t);
    endrule
    rule rule_7668;
        ChannelMessage t;
        t <- mod_5524.get(0);
        mod_4879.put(2, t);
    endrule
    rule rule_7669;
        ChannelMessage t;
        t <- mod_5264.get(0);
        mod_4346.put(2, t);
    endrule
    rule rule_7670;
        ChannelMessage t;
        t <- mod_5462.get(0);
        mod_2378.put(3, t);
    endrule
    rule rule_7671;
        ChannelMessage t;
        t <- mod_5340.get(0);
        mod_3526.put(3, t);
    endrule
    rule rule_7672;
        ChannelMessage t;
        t <- mod_5600.get(75);
        mod_3075.put(1, t);
    endrule
    rule rule_7673;
        ChannelMessage t;
        t <- mod_5491.get(0);
        mod_3649.put(3, t);
    endrule
    rule rule_7674;
        ChannelMessage t;
        t <- mod_5600.get(109);
        mod_4469.put(1, t);
    endrule
    rule rule_7675;
        ChannelMessage t;
        t <- mod_5475.get(0);
        mod_5207.put(3, t);
    endrule
    rule rule_7676;
        ChannelMessage t;
        t <- mod_1189.get(3);
        mod_5443.put(0, t);
    endrule
    rule rule_7677;
        ChannelMessage t;
        t <- mod_4551.get(0);
        mod_5531.put(0, t);
    endrule
    rule rule_7678;
        ChannelMessage t;
        t <- mod_5309.get(123);
        mod_5043.put(0, t);
    endrule
    rule rule_7679;
        ChannelMessage t;
        t <- mod_164.get(3);
        mod_5472.put(0, t);
    endrule
    rule rule_7680;
        ChannelMessage t;
        t <- mod_3075.get(1);
        mod_5466.put(0, t);
    endrule
    rule rule_7681;
        ChannelMessage t;
        t <- mod_164.get(0);
        mod_5489.put(0, t);
    endrule
    rule rule_7682;
        ChannelMessage t;
        t <- mod_779.get(0);
        mod_5639.put(0, t);
    endrule
    rule rule_7683;
        ChannelMessage t;
        t <- mod_1599.get(3);
        mod_5630.put(0, t);
    endrule
    rule rule_7684;
        ChannelMessage t;
        t <- mod_5309.get(124);
        mod_5084.put(0, t);
    endrule
    rule rule_7685;
        ChannelMessage t;
        t <- mod_1476.get(3);
        mod_5313.put(91, t);
    endrule
    rule rule_7686;
        ChannelMessage t;
        t <- mod_2624.get(3);
        mod_5575.put(0, t);
    endrule
    rule rule_7687;
        ChannelMessage t;
        t <- mod_2009.get(0);
        mod_5306.put(0, t);
    endrule
    rule rule_7688;
        ChannelMessage t;
        t <- mod_2829.get(2);
        mod_5591.put(0, t);
    endrule
    rule rule_7689;
        ChannelMessage t;
        t <- mod_5309.get(66);
        mod_2706.put(0, t);
    endrule
    rule rule_7690;
        ChannelMessage t;
        t <- mod_5309.get(126);
        mod_5166.put(0, t);
    endrule
    rule rule_7691;
        ChannelMessage t;
        t <- mod_5448.get(0);
        mod_3198.put(2, t);
    endrule
    rule rule_7692;
        ChannelMessage t;
        t <- mod_5553.get(0);
        mod_3403.put(4, t);
    endrule
    rule rule_7693;
        ChannelMessage t;
        t <- mod_5564.get(0);
        mod_4961.put(2, t);
    endrule
    rule rule_7694;
        ChannelMessage t;
        t <- mod_4428.get(2);
        mod_5250.put(0, t);
    endrule
    rule rule_7695;
        ChannelMessage t;
        t <- mod_1722.get(1);
        mod_5587.put(0, t);
    endrule
    rule rule_7696;
        ChannelMessage t;
        t <- mod_5401.get(0);
        mod_3608.put(4, t);
    endrule
    rule rule_7697;
        ChannelMessage t;
        t <- mod_5635.get(0);
        mod_1558.put(4, t);
    endrule
    rule rule_7698;
        ChannelMessage t;
        t <- mod_2009.get(3);
        mod_5356.put(0, t);
    endrule
    rule rule_7699;
        ChannelMessage t;
        t <- mod_5309.get(13);
        mod_533.put(0, t);
    endrule
    rule rule_7700;
        ChannelMessage t;
        t <- mod_1230.get(2);
        mod_5530.put(0, t);
    endrule
    rule rule_7701;
        ChannelMessage t;
        t <- mod_5600.get(90);
        mod_3690.put(1, t);
    endrule
    rule rule_7702;
        ChannelMessage t;
        t <- mod_2542.get(0);
        mod_5429.put(0, t);
    endrule
    rule rule_7703;
        ChannelMessage t;
        t <- mod_4879.get(0);
        mod_5613.put(0, t);
    endrule
    rule rule_7704;
        ChannelMessage t;
        t <- mod_3485.get(0);
        mod_5588.put(0, t);
    endrule
    rule rule_7705;
        ChannelMessage t;
        t <- mod_5309.get(117);
        mod_4797.put(0, t);
    endrule
    rule rule_7706;
        ChannelMessage t;
        t <- mod_5640.get(0);
        mod_5166.put(3, t);
    endrule
    rule rule_7707;
        ChannelMessage t;
        t <- mod_4920.get(2);
        mod_5294.put(0, t);
    endrule
    rule rule_7708;
        ChannelMessage t;
        t <- mod_1722.get(3);
        mod_5450.put(0, t);
    endrule
    rule rule_7709;
        ChannelMessage t;
        t <- mod_5405.get(0);
        mod_820.put(3, t);
    endrule
    rule rule_7710;
        ChannelMessage t;
        t <- mod_1066.get(0);
        mod_5313.put(101, t);
    endrule
    rule rule_7711;
        ChannelMessage t;
        t <- mod_5600.get(93);
        mod_3813.put(1, t);
    endrule
    rule rule_7712;
        ChannelMessage t;
        t <- mod_5387.get(0);
        mod_1189.put(3, t);
    endrule
    rule rule_7713;
        ChannelMessage t;
        t <- mod_5445.get(0);
        mod_82.put(2, t);
    endrule
    rule rule_7714;
        ChannelMessage t;
        t <- mod_1476.get(1);
        mod_5617.put(0, t);
    endrule
    rule rule_7715;
        ChannelMessage t;
        t <- mod_5600.get(115);
        mod_4715.put(1, t);
    endrule
    rule rule_7716;
        ChannelMessage t;
        t <- mod_5337.get(0);
        mod_246.put(2, t);
    endrule
    rule rule_7717;
        ChannelMessage t;
        t <- mod_5600.get(20);
        mod_820.put(1, t);
    endrule
    rule rule_7718;
        ChannelMessage t;
        t <- mod_5514.get(0);
        mod_2952.put(4, t);
    endrule
    rule rule_7719;
        ChannelMessage t;
        t <- mod_5309.get(52);
        mod_2132.put(0, t);
    endrule
    rule rule_7720;
        ChannelMessage t;
        t <- mod_4059.get(2);
        mod_5366.put(0, t);
    endrule
    rule rule_7721;
        ChannelMessage t;
        t <- mod_5525.get(0);
        mod_4387.put(4, t);
    endrule
    rule rule_7722;
        ChannelMessage t;
        t <- mod_5385.get(0);
        mod_574.put(4, t);
    endrule
    rule rule_7723;
        ChannelMessage t;
        t <- mod_5600.get(99);
        mod_4059.put(1, t);
    endrule
    rule rule_7724;
        ChannelMessage t;
        t <- mod_1886.get(0);
        mod_5602.put(0, t);
    endrule
    rule rule_7725;
        ChannelMessage t;
        t <- mod_5429.get(0);
        mod_2542.put(2, t);
    endrule
    rule rule_7726;
        ChannelMessage t;
        t <- mod_5309.get(70);
        mod_2870.put(0, t);
    endrule
    rule rule_7727;
        ChannelMessage t;
        t <- mod_5440.get(0);
        mod_1886.put(4, t);
    endrule
    rule rule_7728;
        ChannelMessage t;
        t <- mod_5581.get(0);
        mod_1476.put(4, t);
    endrule
    rule rule_7729;
        ChannelMessage t;
        t <- mod_5309.get(81);
        mod_3321.put(0, t);
    endrule
    rule rule_7730;
        ChannelMessage t;
        t <- mod_2665.get(0);
        mod_5595.put(0, t);
    endrule
    rule rule_7731;
        ChannelMessage t;
        t <- mod_5549.get(0);
        mod_861.put(2, t);
    endrule
    rule rule_7732;
        ChannelMessage t;
        t <- mod_5309.get(82);
        mod_3362.put(0, t);
    endrule
    rule rule_7733;
        ChannelMessage t;
        t <- mod_5600.get(100);
        mod_4100.put(1, t);
    endrule
    rule rule_7734;
        ChannelMessage t;
        t <- mod_820.get(3);
        mod_5313.put(107, t);
    endrule
    rule rule_7735;
        ChannelMessage t;
        t <- mod_5357.get(0);
        mod_4961.put(3, t);
    endrule
    rule rule_7736;
        ChannelMessage t;
        t <- mod_5620.get(0);
        mod_5002.put(4, t);
    endrule
    rule rule_7737;
        ChannelMessage t;
        t <- mod_5600.get(35);
        mod_1435.put(1, t);
    endrule
    rule rule_7738;
        ChannelMessage t;
        t <- mod_5309.get(3);
        mod_123.put(0, t);
    endrule
    rule rule_7739;
        ChannelMessage t;
        t <- mod_5600.get(32);
        mod_1312.put(1, t);
    endrule
    rule rule_7740;
        ChannelMessage t;
        t <- mod_1517.get(3);
        mod_5313.put(90, t);
    endrule
    rule rule_7741;
        ChannelMessage t;
        t <- mod_2952.get(0);
        mod_5378.put(0, t);
    endrule
    rule rule_7742;
        ChannelMessage t;
        t <- mod_4592.get(3);
        mod_5442.put(0, t);
    endrule
    rule rule_7743;
        ChannelMessage t;
        t <- mod_5546.get(0);
        mod_5125.put(2, t);
    endrule
    rule rule_7744;
        ChannelMessage t;
        t <- mod_5600.get(18);
        mod_738.put(1, t);
    endrule
    rule rule_7745;
        ChannelMessage t;
        t <- mod_4346.get(3);
        mod_5313.put(21, t);
    endrule
    rule rule_7746;
        ChannelMessage t;
        t <- mod_5600.get(67);
        mod_2747.put(1, t);
    endrule
    rule rule_7747;
        ChannelMessage t;
        t <- mod_2870.get(3);
        mod_5454.put(0, t);
    endrule
    rule rule_7748;
        ChannelMessage t;
        t <- mod_5518.get(0);
        mod_2911.put(2, t);
    endrule
    rule rule_7749;
        ChannelMessage t;
        t <- mod_5473.get(0);
        mod_451.put(4, t);
    endrule
    rule rule_7750;
        ChannelMessage t;
        t <- mod_3731.get(2);
        mod_5496.put(0, t);
    endrule
    rule rule_7751;
        ChannelMessage t;
        t <- mod_4838.get(3);
        mod_5598.put(0, t);
    endrule
    rule rule_7752;
        ChannelMessage t;
        t <- mod_5447.get(0);
        mod_3362.put(2, t);
    endrule
    rule rule_7753;
        ChannelMessage t;
        t <- mod_4100.get(0);
        mod_5499.put(0, t);
    endrule
    rule rule_7754;
        ChannelMessage t;
        t <- mod_4428.get(0);
        mod_5627.put(0, t);
    endrule
    rule rule_7755;
        ChannelMessage t;
        t <- mod_2132.get(1);
        mod_5291.put(0, t);
    endrule
    rule rule_7756;
        ChannelMessage t;
        t <- mod_3731.get(0);
        mod_5642.put(0, t);
    endrule
    rule rule_7757;
        ChannelMessage t;
        t <- mod_5260.get(0);
        mod_1148.put(3, t);
    endrule
    rule rule_7758;
        ChannelMessage t;
        t <- mod_2091.get(2);
        mod_5313.put(76, t);
    endrule
    rule rule_7759;
        ChannelMessage t;
        t <- mod_3075.get(0);
        mod_5464.put(0, t);
    endrule
    rule rule_7760;
        ChannelMessage t;
        t <- mod_5309.get(60);
        mod_2460.put(0, t);
    endrule
    rule rule_7761;
        ChannelMessage t;
        t <- mod_5323.get(0);
        mod_3362.put(3, t);
    endrule
    rule rule_7762;
        ChannelMessage t;
        t <- mod_902.get(3);
        mod_5547.put(0, t);
    endrule
    rule rule_7763;
        ChannelMessage t;
        t <- mod_5263.get(0);
        mod_4387.put(3, t);
    endrule
    rule rule_7764;
        ChannelMessage t;
        t <- mod_1681.get(2);
        mod_5313.put(86, t);
    endrule
    rule rule_7765;
        ChannelMessage t;
        t <- mod_5309.get(39);
        mod_1599.put(0, t);
    endrule
    rule rule_7766;
        ChannelMessage t;
        t <- mod_5309.get(46);
        mod_1886.put(0, t);
    endrule
    rule rule_7767;
        ChannelMessage t;
        t <- mod_5336.get(0);
        mod_4264.put(4, t);
    endrule
    rule rule_7768;
        ChannelMessage t;
        t <- mod_5125.get(2);
        mod_5546.put(0, t);
    endrule
    rule rule_7769;
        ChannelMessage t;
        t <- mod_5420.get(0);
        mod_2214.put(4, t);
    endrule
    rule rule_7770;
        ChannelMessage t;
        t <- mod_861.get(3);
        mod_5549.put(0, t);
    endrule
    rule rule_7771;
        ChannelMessage t;
        t <- mod_5309.get(76);
        mod_3116.put(0, t);
    endrule
    rule rule_7772;
        ChannelMessage t;
        t <- mod_5468.get(0);
        mod_4100.put(4, t);
    endrule
    rule rule_7773;
        ChannelMessage t;
        t <- mod_5578.get(0);
        mod_1599.put(2, t);
    endrule
    rule rule_7774;
        ChannelMessage t;
        t <- mod_5322.get(0);
        mod_3854.put(4, t);
    endrule
    rule rule_7775;
        ChannelMessage t;
        t <- mod_5502.get(0);
        mod_2337.put(2, t);
    endrule
    rule rule_7776;
        ChannelMessage t;
        t <- mod_4059.get(3);
        mod_5560.put(0, t);
    endrule
    rule rule_7777;
        ChannelMessage t;
        t <- mod_943.get(3);
        mod_5313.put(104, t);
    endrule
    rule rule_7778;
        ChannelMessage t;
        t <- mod_123.get(1);
        mod_5313.put(124, t);
    endrule
    rule rule_7779;
        ChannelMessage t;
        t <- mod_3198.get(3);
        mod_5507.put(0, t);
    endrule
    rule rule_7780;
        ChannelMessage t;
        t <- mod_5284.get(0);
        mod_1353.put(3, t);
    endrule
    rule rule_7781;
        ChannelMessage t;
        t <- mod_5509.get(0);
        mod_4510.put(2, t);
    endrule
    rule rule_7782;
        ChannelMessage t;
        t <- mod_4100.get(2);
        mod_5468.put(0, t);
    endrule
    rule rule_7783;
        ChannelMessage t;
        t <- mod_3854.get(1);
        mod_5593.put(0, t);
    endrule
    rule rule_7784;
        ChannelMessage t;
        t <- mod_5301.get(0);
        mod_1271.put(4, t);
    endrule
    rule rule_7785;
        ChannelMessage t;
        t <- mod_5600.get(55);
        mod_2255.put(1, t);
    endrule
    rule rule_7786;
        ChannelMessage t;
        t <- mod_5600.get(91);
        mod_3731.put(1, t);
    endrule
    rule rule_7787;
        ChannelMessage t;
        t <- mod_574.get(2);
        mod_5455.put(0, t);
    endrule
    rule rule_7788;
        ChannelMessage t;
        t <- mod_3895.get(3);
        mod_5544.put(0, t);
    endrule
    rule rule_7789;
        ChannelMessage t;
        t <- mod_5306.get(0);
        mod_2009.put(3, t);
    endrule
    rule rule_7790;
        ChannelMessage t;
        t <- mod_5327.get(0);
        mod_4182.put(3, t);
    endrule
    rule rule_7791;
        ChannelMessage t;
        t <- mod_2788.get(0);
        mod_5645.put(0, t);
    endrule
    rule rule_7792;
        ChannelMessage t;
        t <- mod_5643.get(0);
        mod_4223.put(4, t);
    endrule
    rule rule_7793;
        ChannelMessage t;
        t <- mod_5464.get(0);
        mod_3075.put(2, t);
    endrule
    rule rule_7794;
        ChannelMessage t;
        t <- mod_5470.get(0);
        mod_3116.put(4, t);
    endrule
    rule rule_7795;
        ChannelMessage t;
        t <- mod_5422.get(0);
        mod_2747.put(2, t);
    endrule
    rule rule_7796;
        ChannelMessage t;
        t <- mod_5444.get(0);
        mod_2419.put(2, t);
    endrule
    rule rule_7797;
        ChannelMessage t;
        t <- mod_5310.get(0);
        mod_1927.put(4, t);
    endrule
    rule rule_7798;
        ChannelMessage t;
        t <- mod_2460.get(1);
        mod_5313.put(67, t);
    endrule
    rule rule_7799;
        ChannelMessage t;
        t <- mod_41.get(3);
        mod_5570.put(0, t);
    endrule
    rule rule_7800;
        ChannelMessage t;
        t <- mod_5287.get(0);
        mod_2829.put(2, t);
    endrule
    rule rule_7801;
        ChannelMessage t;
        t <- mod_5309.get(41);
        mod_1681.put(0, t);
    endrule
    rule rule_7802;
        ChannelMessage t;
        t <- mod_5600.get(101);
        mod_4141.put(1, t);
    endrule
    rule rule_7803;
        ChannelMessage t;
        t <- mod_5283.get(0);
        mod_1435.put(3, t);
    endrule
    rule rule_7804;
        ChannelMessage t;
        t <- mod_5304.get(0);
        mod_1312.put(2, t);
    endrule
    rule rule_7805;
        ChannelMessage t;
        t <- mod_5274.get(0);
        mod_5043.put(4, t);
    endrule
    rule rule_7806;
        ChannelMessage t;
        t <- mod_5413.get(0);
        mod_4305.put(2, t);
    endrule
    rule rule_7807;
        ChannelMessage t;
        t <- mod_533.get(1);
        mod_5316.put(0, t);
    endrule
    rule rule_7808;
        ChannelMessage t;
        t <- mod_2460.get(2);
        mod_5338.put(0, t);
    endrule
    rule rule_7809;
        ChannelMessage t;
        t <- mod_4633.get(3);
        mod_5532.put(0, t);
    endrule
    rule rule_7810;
        ChannelMessage t;
        t <- mod_5002.get(2);
        mod_5620.put(0, t);
    endrule
    rule rule_7811;
        ChannelMessage t;
        t <- mod_2542.get(1);
        mod_5286.put(0, t);
    endrule
    rule rule_7812;
        ChannelMessage t;
        t <- mod_3444.get(0);
        mod_5384.put(0, t);
    endrule
    rule rule_7813;
        ChannelMessage t;
        t <- mod_5280.get(0);
        mod_3936.put(3, t);
    endrule
    rule rule_7814;
        ChannelMessage t;
        t <- mod_5551.get(0);
        mod_2296.put(4, t);
    endrule
    rule rule_7815;
        ChannelMessage t;
        t <- mod_5600.get(1);
        mod_41.put(1, t);
    endrule
    rule rule_7816;
        ChannelMessage t;
        t <- mod_5531.get(0);
        mod_4551.put(3, t);
    endrule
    rule rule_7817;
        ChannelMessage t;
        t <- mod_5600.get(26);
        mod_1066.put(1, t);
    endrule
    rule rule_7818;
        ChannelMessage t;
        t <- mod_5609.get(0);
        mod_4182.put(2, t);
    endrule
    rule rule_7819;
        ChannelMessage t;
        t <- mod_738.get(0);
        mod_5381.put(0, t);
    endrule
    rule rule_7820;
        ChannelMessage t;
        t <- mod_1558.get(0);
        mod_5635.put(0, t);
    endrule
    rule rule_7821;
        ChannelMessage t;
        t <- mod_2911.get(0);
        mod_5313.put(56, t);
    endrule
    rule rule_7822;
        ChannelMessage t;
        t <- mod_3936.get(1);
        mod_5476.put(0, t);
    endrule
    rule rule_7823;
        ChannelMessage t;
        t <- mod_3239.get(3);
        mod_5342.put(0, t);
    endrule
    rule rule_7824;
        ChannelMessage t;
        t <- mod_5403.get(0);
        mod_2091.put(2, t);
    endrule
    rule rule_7825;
        ChannelMessage t;
        t <- mod_5309.get(113);
        mod_4633.put(0, t);
    endrule
    rule rule_7826;
        ChannelMessage t;
        t <- mod_2747.get(3);
        mod_5485.put(0, t);
    endrule
    rule rule_7827;
        ChannelMessage t;
        t <- mod_5266.get(0);
        mod_3157.put(3, t);
    endrule
    rule rule_7828;
        ChannelMessage t;
        t <- mod_5309.get(99);
        mod_4059.put(0, t);
    endrule
    rule rule_7829;
        ChannelMessage t;
        t <- mod_5309.get(125);
        mod_5125.put(0, t);
    endrule
    rule rule_7830;
        ChannelMessage t;
        t <- mod_5583.get(0);
        mod_1189.put(4, t);
    endrule
    rule rule_7831;
        ChannelMessage t;
        t <- mod_5257.get(0);
        mod_1599.put(4, t);
    endrule
    rule rule_7832;
        ChannelMessage t;
        t <- mod_5277.get(0);
        mod_1804.put(3, t);
    endrule
    rule rule_7833;
        ChannelMessage t;
        t <- mod_1681.get(3);
        mod_5312.put(0, t);
    endrule
    rule rule_7834;
        ChannelMessage t;
        t <- mod_328.get(1);
        mod_5251.put(0, t);
    endrule
    rule rule_7835;
        ChannelMessage t;
        t <- mod_5622.get(0);
        mod_4879.put(4, t);
    endrule
    rule rule_7836;
        ChannelMessage t;
        t <- mod_3977.get(3);
        mod_5493.put(0, t);
    endrule
    rule rule_7837;
        ChannelMessage t;
        t <- mod_5460.get(0);
        mod_5600.put(0, t);
    endrule
    rule rule_7838;
        ChannelMessage t;
        t <- mod_5621.get(0);
        mod_2911.put(3, t);
    endrule
    rule rule_7839;
        ChannelMessage t;
        t <- mod_5309.get(106);
        mod_4346.put(0, t);
    endrule
    rule rule_7840;
        ChannelMessage t;
        t <- mod_5374.get(0);
        mod_2665.put(3, t);
    endrule
    rule rule_7841;
        ChannelMessage t;
        t <- mod_4510.get(1);
        mod_5368.put(0, t);
    endrule
    rule rule_7842;
        ChannelMessage t;
        t <- mod_574.get(1);
        mod_5313.put(113, t);
    endrule
    rule rule_7843;
        ChannelMessage t;
        t <- mod_943.get(2);
        mod_5490.put(0, t);
    endrule
    rule rule_7844;
        ChannelMessage t;
        t <- mod_5600.get(117);
        mod_4797.put(1, t);
    endrule
    rule rule_7845;
        ChannelMessage t;
        t <- mod_697.get(1);
        mod_5298.put(0, t);
    endrule
    rule rule_7846;
        ChannelMessage t;
        t <- mod_1025.get(1);
        mod_5423.put(0, t);
    endrule
    rule rule_7847;
        ChannelMessage t;
        t <- mod_5309.get(87);
        mod_3567.put(0, t);
    endrule
    rule rule_7848;
        ChannelMessage t;
        t <- mod_41.get(2);
        mod_5313.put(126, t);
    endrule
    rule rule_7849;
        ChannelMessage t;
        t <- mod_5342.get(0);
        mod_3239.put(3, t);
    endrule
    rule rule_7850;
        ChannelMessage t;
        t <- mod_5309.get(112);
        mod_4592.put(0, t);
    endrule
    rule rule_7851;
        ChannelMessage t;
        t <- mod_1886.get(1);
        mod_5440.put(0, t);
    endrule
    rule rule_7852;
        ChannelMessage t;
        t <- mod_5600.get(17);
        mod_697.put(1, t);
    endrule
    rule rule_7853;
        ChannelMessage t;
        t <- mod_2624.get(1);
        mod_5313.put(63, t);
    endrule
    rule rule_7854;
        ChannelMessage t;
        t <- mod_5618.get(0);
        mod_3485.put(4, t);
    endrule
    rule rule_7855;
        ChannelMessage t;
        t <- mod_3157.get(3);
        mod_5355.put(0, t);
    endrule
    rule rule_7856;
        ChannelMessage t;
        t <- mod_2911.get(1);
        mod_5621.put(0, t);
    endrule
    rule rule_7857;
        ChannelMessage t;
        t <- mod_5267.get(0);
        mod_410.put(3, t);
    endrule
    rule rule_7858;
        ChannelMessage t;
        t <- mod_5501.get(0);
        mod_3649.put(4, t);
    endrule
    rule rule_7859;
        ChannelMessage t;
        t <- mod_5600.get(107);
        mod_4387.put(1, t);
    endrule
    rule rule_7860;
        ChannelMessage t;
        t <- mod_5590.get(0);
        mod_2214.put(2, t);
    endrule
    rule rule_7861;
        ChannelMessage t;
        t <- mod_3362.get(3);
        mod_5302.put(0, t);
    endrule
    rule rule_7862;
        ChannelMessage t;
        t <- mod_2132.get(3);
        mod_5313.put(75, t);
    endrule
    rule rule_7863;
        ChannelMessage t;
        t <- mod_5588.get(0);
        mod_3485.put(2, t);
    endrule
    rule rule_7864;
        ChannelMessage t;
        t <- mod_4715.get(3);
        mod_5567.put(0, t);
    endrule
    rule rule_7865;
        ChannelMessage t;
        t <- mod_1394.get(3);
        mod_5592.put(0, t);
    endrule
    rule rule_7866;
        ChannelMessage t;
        t <- mod_5398.get(0);
        mod_3567.put(2, t);
    endrule
    rule rule_7867;
        ChannelMessage t;
        t <- mod_5600.get(72);
        mod_2952.put(1, t);
    endrule
    rule rule_7868;
        ChannelMessage t;
        t <- mod_123.get(0);
        mod_5328.put(0, t);
    endrule
    rule rule_7869;
        ChannelMessage t;
        t <- mod_5636.get(0);
        mod_3034.put(4, t);
    endrule
    rule rule_7870;
        ChannelMessage t;
        t <- mod_5600.get(104);
        mod_4264.put(1, t);
    endrule
    rule rule_7871;
        ChannelMessage t;
        t <- mod_1886.get(3);
        mod_5542.put(0, t);
    endrule
    rule rule_7872;
        ChannelMessage t;
        t <- mod_4715.get(0);
        mod_5373.put(0, t);
    endrule
    rule rule_7873;
        ChannelMessage t;
        t <- mod_4674.get(3);
        mod_5375.put(0, t);
    endrule
    rule rule_7874;
        ChannelMessage t;
        t <- mod_5523.get(0);
        mod_5313.put(128, t);
    endrule
    rule rule_7875;
        ChannelMessage t;
        t <- mod_5343.get(0);
        mod_615.put(4, t);
    endrule
    rule rule_7876;
        ChannelMessage t;
        t <- mod_3526.get(2);
        mod_5340.put(0, t);
    endrule
    rule rule_7877;
        ChannelMessage t;
        t <- mod_3034.get(1);
        mod_5252.put(0, t);
    endrule
    rule rule_7878;
        ChannelMessage t;
        t <- mod_5309.get(1);
        mod_41.put(0, t);
    endrule
    rule rule_7879;
        ChannelMessage t;
        t <- mod_5600.get(69);
        mod_2829.put(1, t);
    endrule
    rule rule_7880;
        ChannelMessage t;
        t <- mod_5372.get(1);
        mod_5495.put(0, t);
    endrule
    rule rule_7881;
        ChannelMessage t;
        t <- mod_5573.get(0);
        mod_2173.put(3, t);
    endrule
    rule rule_7882;
        ChannelMessage t;
        t <- mod_4633.get(1);
        mod_5313.put(14, t);
    endrule
    rule rule_7883;
        ChannelMessage t;
        t <- mod_4469.get(2);
        mod_5313.put(18, t);
    endrule
    rule rule_7884;
        ChannelMessage t;
        t <- mod_5289.get(0);
        mod_4018.put(4, t);
    endrule
    rule rule_7885;
        ChannelMessage t;
        t <- mod_5309.get(73);
        mod_2993.put(0, t);
    endrule
    rule rule_7886;
        ChannelMessage t;
        t <- mod_5406.get(0);
        mod_2706.put(4, t);
    endrule
    rule rule_7887;
        ChannelMessage t;
        t <- mod_5597.get(0);
        mod_1148.put(4, t);
    endrule
    rule rule_7888;
        ChannelMessage t;
        t <- mod_5043.get(3);
        mod_5313.put(4, t);
    endrule
    rule rule_7889;
        ChannelMessage t;
        t <- mod_4510.get(0);
        mod_5313.put(17, t);
    endrule
    rule rule_7890;
        ChannelMessage t;
        t <- mod_3157.get(0);
        mod_5647.put(0, t);
    endrule
    rule rule_7891;
        ChannelMessage t;
        t <- mod_5207.get(0);
        mod_5313.put(0, t);
    endrule
    rule rule_7892;
        ChannelMessage t;
        t <- mod_5600.get(47);
        mod_1927.put(1, t);
    endrule
    rule rule_7893;
        ChannelMessage t;
        t <- mod_3690.get(0);
        mod_5607.put(0, t);
    endrule
    rule rule_7894;
        ChannelMessage t;
        t <- mod_1025.get(3);
        mod_5313.put(102, t);
    endrule
    rule rule_7895;
        ChannelMessage t;
        t <- mod_5570.get(0);
        mod_41.put(4, t);
    endrule
    rule rule_7896;
        ChannelMessage t;
        t <- mod_5309.get(24);
        mod_984.put(0, t);
    endrule
    rule rule_7897;
        ChannelMessage t;
        t <- mod_1435.get(3);
        mod_5313.put(92, t);
    endrule
    rule rule_7898;
        ChannelMessage t;
        t <- mod_5002.get(1);
        mod_5388.put(0, t);
    endrule
    rule rule_7899;
        ChannelMessage t;
        t <- mod_5309.get(48);
        mod_1968.put(0, t);
    endrule
    rule rule_7900;
        ChannelMessage t;
        t <- mod_5309.get(100);
        mod_4100.put(0, t);
    endrule
    rule rule_7901;
        ChannelMessage t;
        t <- mod_5600.get(81);
        mod_3321.put(1, t);
    endrule
    rule rule_7902;
        ChannelMessage t;
        t <- mod_2706.get(2);
        mod_5297.put(0, t);
    endrule
    rule rule_7903;
        ChannelMessage t;
        t <- mod_4141.get(1);
        mod_5410.put(0, t);
    endrule
    rule rule_7904;
        ChannelMessage t;
        t <- mod_3075.get(3);
        mod_5313.put(52, t);
    endrule
    rule rule_7905;
        ChannelMessage t;
        t <- mod_4674.get(0);
        mod_5634.put(0, t);
    endrule
    rule rule_7906;
        ChannelMessage t;
        t <- mod_3157.get(2);
        mod_5313.put(50, t);
    endrule
    rule rule_7907;
        ChannelMessage t;
        t <- mod_1066.get(2);
        mod_5308.put(0, t);
    endrule
    rule rule_7908;
        ChannelMessage t;
        t <- mod_2870.get(1);
        mod_5629.put(0, t);
    endrule
    rule rule_7909;
        ChannelMessage t;
        t <- mod_1804.get(1);
        mod_5313.put(83, t);
    endrule
    rule rule_7910;
        ChannelMessage t;
        t <- mod_5365.get(0);
        mod_2378.put(4, t);
    endrule
    rule rule_7911;
        ChannelMessage t;
        t <- mod_5397.get(0);
        mod_4838.put(4, t);
    endrule
    rule rule_7912;
        ChannelMessage t;
        t <- mod_5481.get(0);
        mod_5526.put(0, t);
    endrule
    rule rule_7913;
        ChannelMessage t;
        t <- mod_5511.get(0);
        mod_4223.put(3, t);
    endrule
    rule rule_7914;
        ChannelMessage t;
        t <- mod_861.get(1);
        mod_5285.put(0, t);
    endrule
    rule rule_7915;
        ChannelMessage t;
        t <- mod_1353.get(0);
        mod_5284.put(0, t);
    endrule
    rule rule_7916;
        ChannelMessage t;
        t <- mod_3362.get(1);
        mod_5447.put(0, t);
    endrule
    rule rule_7917;
        ChannelMessage t;
        t <- mod_5600.get(97);
        mod_3977.put(1, t);
    endrule
    rule rule_7918;
        ChannelMessage t;
        t <- mod_5600.get(124);
        mod_5084.put(1, t);
    endrule
    rule rule_7919;
        ChannelMessage t;
        t <- mod_3936.get(0);
        mod_5256.put(0, t);
    endrule
    rule rule_7920;
        ChannelMessage t;
        t <- mod_3567.get(2);
        mod_5398.put(0, t);
    endrule
    rule rule_7921;
        ChannelMessage t;
        t <- mod_5312.get(0);
        mod_1681.put(3, t);
    endrule
    rule rule_7922;
        ChannelMessage t;
        t <- mod_3731.get(1);
        mod_5487.put(0, t);
    endrule
    rule rule_7923;
        ChannelMessage t;
        t <- mod_5309.get(50);
        mod_2050.put(0, t);
    endrule
    rule rule_7924;
        ChannelMessage t;
        t <- mod_5317.get(0);
        mod_4715.put(3, t);
    endrule
    rule rule_7925;
        ChannelMessage t;
        t <- mod_5307.get(0);
        mod_738.put(4, t);
    endrule
    rule rule_7926;
        ChannelMessage t;
        t <- mod_5084.get(1);
        mod_5418.put(0, t);
    endrule
    rule rule_7927;
        ChannelMessage t;
        t <- mod_5309.get(78);
        mod_3198.put(0, t);
    endrule
    rule rule_7928;
        ChannelMessage t;
        t <- mod_5309.get(54);
        mod_2214.put(0, t);
    endrule
    rule rule_7929;
        ChannelMessage t;
        t <- mod_5383.get(0);
        mod_3198.put(4, t);
    endrule
    rule rule_7930;
        ChannelMessage t;
        t <- mod_410.get(1);
        mod_5399.put(0, t);
    endrule
    rule rule_7931;
        ChannelMessage t;
        t <- mod_2337.get(2);
        mod_5522.put(0, t);
    endrule
    rule rule_7932;
        ChannelMessage t;
        t <- mod_3772.get(0);
        mod_5279.put(0, t);
    endrule
    rule rule_7933;
        ChannelMessage t;
        t <- mod_5538.get(0);
        mod_1968.put(3, t);
    endrule
    rule rule_7934;
        ChannelMessage t;
        t <- mod_5600.get(15);
        mod_615.put(1, t);
    endrule
    rule rule_7935;
        ChannelMessage t;
        t <- mod_5309.get(15);
        mod_615.put(0, t);
    endrule
    rule rule_7936;
        ChannelMessage t;
        t <- mod_5600.get(57);
        mod_2337.put(1, t);
    endrule
    rule rule_7937;
        ChannelMessage t;
        t <- mod_5598.get(0);
        mod_4838.put(2, t);
    endrule
    rule rule_7938;
        ChannelMessage t;
        t <- mod_1763.get(3);
        mod_5409.put(0, t);
    endrule
    rule rule_7939;
        ChannelMessage t;
        t <- mod_1763.get(2);
        mod_5290.put(0, t);
    endrule
    rule rule_7940;
        ChannelMessage t;
        t <- mod_5552.get(0);
        mod_5002.put(3, t);
    endrule
    rule rule_7941;
        ChannelMessage t;
        t <- mod_615.get(3);
        mod_5474.put(0, t);
    endrule
    rule rule_7942;
        ChannelMessage t;
        t <- mod_5446.get(0);
        mod_5125.put(4, t);
    endrule
    rule rule_7943;
        ChannelMessage t;
        t <- mod_5566.get(0);
        mod_164.put(3, t);
    endrule
    rule rule_7944;
        ChannelMessage t;
        t <- mod_1558.get(2);
        mod_5269.put(0, t);
    endrule
    rule rule_7945;
        ChannelMessage t;
        t <- mod_4756.get(1);
        mod_5278.put(0, t);
    endrule
    rule rule_7946;
        ChannelMessage t;
        t <- mod_5321.get(0);
        mod_2009.put(4, t);
    endrule
    rule rule_7947;
        ChannelMessage t;
        t <- mod_5384.get(0);
        mod_3444.put(4, t);
    endrule
    rule rule_7948;
        ChannelMessage t;
        t <- mod_5399.get(0);
        mod_410.put(4, t);
    endrule
    rule rule_7949;
        ChannelMessage t;
        t <- mod_5412.get(0);
        mod_2993.put(2, t);
    endrule
    rule rule_7950;
        ChannelMessage t;
        t <- mod_779.get(3);
        mod_5313.put(108, t);
    endrule
    rule rule_7951;
        ChannelMessage t;
        t <- mod_2501.get(3);
        mod_5363.put(0, t);
    endrule
    rule rule_7952;
        ChannelMessage t;
        t <- mod_3116.get(3);
        mod_5543.put(0, t);
    endrule

endmodule
endpackage
