package Step;
import Operation::*;
import Types::*;
import Vector::*;
import FShow::*;
import Debug::*;
import PMU::*;
import RamulatorArbiter::*;
import RandomLoad::*;

(* synthesize *)
module mkHypernode (Operation_IFC);
    Operation_IFC mod_1_inner <- mkReshape(2, 64);
    Operation_IFC mod_1 <- mkDebugOperation(mod_1_inner, "mod_1");
    Operation_IFC mod_2_inner <- mkFlatten(1);
    Operation_IFC mod_2 <- mkDebugOperation(mod_2_inner, "mod_2");
    Operation_IFC mod_3_inner <- mkFlatten(2);
    Operation_IFC mod_3 <- mkDebugOperation(mod_3_inner, "mod_3");
    Operation_IFC mod_4_inner <- mkAccumBigTile(retile_row_tile, 3);
    Operation_IFC mod_4 <- mkDebugOperation(mod_4_inner, "mod_4");
    Broadcast_IFC#(4) mod_5_inner <- mkBroadcast(4);
    Operation_IFC mod_5 <- mkDebugOperation(mod_5_inner.op, "mod_5");
    PMU_IFC mod_6_bufferize <- mkPMU(2);
    Operation_IFC mod_6_inner = mod_6_bufferize.operation;
    Operation_IFC mod_6 <- mkDebugOperation(mod_6_inner, "mod_6");
    Broadcast_IFC#(2) mod_7_inner <- mkBroadcast(2);
    Operation_IFC mod_7 <- mkDebugOperation(mod_7_inner.op, "mod_7");
    PMU_IFC mod_8_bufferize <- mkPMU(1);
    Operation_IFC mod_8_inner = mod_8_bufferize.operation;
    Operation_IFC mod_8 <- mkDebugOperation(mod_8_inner, "mod_8");
    Operation_IFC mod_9_inner <- mkBinaryMap(1156, matmul_t_tile);
    Operation_IFC mod_9 <- mkDebugOperation(mod_9_inner, "mod_9");
    Operation_IFC mod_10_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_10 <- mkDebugOperation(mod_10_inner, "mod_10");
    Operation_IFC mod_11_inner <- mkBinaryMap(1924, mul_tile);
    Operation_IFC mod_11 <- mkDebugOperation(mod_11_inner, "mod_11");
    PMU_IFC mod_12_bufferize <- mkPMU(1);
    Operation_IFC mod_12_inner = mod_12_bufferize.operation;
    Operation_IFC mod_12 <- mkDebugOperation(mod_12_inner, "mod_12");
    Operation_IFC mod_13_inner <- mkBinaryMap(2563, matmul_t_tile);
    Operation_IFC mod_13 <- mkDebugOperation(mod_13_inner, "mod_13");
    Operation_IFC mod_14_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_14 <- mkDebugOperation(mod_14_inner, "mod_14");
    Operation_IFC mod_15_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_15 <- mkDebugOperation(mod_15_inner, "mod_15");
    Operation_IFC mod_16_inner <- mkTiledRetileStreamify(3, True, True);
    Operation_IFC mod_16 <- mkDebugOperation(mod_16_inner, "mod_16");
    Operation_IFC mod_17_inner <- mkBinaryMap(2823, mul_tile);
    Operation_IFC mod_17 <- mkDebugOperation(mod_17_inner, "mod_17");
    PMU_IFC mod_18_bufferize <- mkPMU(1);
    Operation_IFC mod_18_inner = mod_18_bufferize.operation;
    Operation_IFC mod_18 <- mkDebugOperation(mod_18_inner, "mod_18");
    PMU_IFC mod_19_bufferize <- mkPMU(2);
    Operation_IFC mod_19_inner = mod_19_bufferize.operation;
    Operation_IFC mod_19 <- mkDebugOperation(mod_19_inner, "mod_19");
    PMU_IFC mod_20_bufferize <- mkPMU(2);
    Operation_IFC mod_20_inner = mod_20_bufferize.operation;
    Operation_IFC mod_20 <- mkDebugOperation(mod_20_inner, "mod_20");
    Operation_IFC mod_21_inner <- mkRepeatStatic(8);
    Operation_IFC mod_21 <- mkDebugOperation(mod_21_inner, "mod_21");
    Operation_IFC mod_22_inner <- mkFlatten(1);
    Operation_IFC mod_22 <- mkDebugOperation(mod_22_inner, "mod_22");
    Operation_IFC mod_23_inner <- mkFlatten(0);
    Operation_IFC mod_23 <- mkDebugOperation(mod_23_inner, "mod_23");
    Operation_IFC mod_24_inner <- mkDynamicRandomLoad(Cons(1, Cons(2, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_24 <- mkDebugOperation(mod_24_inner, "mod_24");
    Operation_IFC mod_25_inner <- mkRepeatStatic(3);
    Operation_IFC mod_25 <- mkDebugOperation(mod_25_inner, "mod_25");
    Operation_IFC mod_26_inner <- mkUnaryMap(1796, silu_tile);
    Operation_IFC mod_26 <- mkDebugOperation(mod_26_inner, "mod_26");
    Operation_IFC mod_27_inner <- mkAccum(add_tile, 1);
    Operation_IFC mod_27 <- mkDebugOperation(mod_27_inner, "mod_27");
    Operation_IFC mod_28_inner <- mkBinaryMap(1668, matmul_t_tile);
    Operation_IFC mod_28 <- mkDebugOperation(mod_28_inner, "mod_28");
    PMU_IFC mod_29_bufferize <- mkPMU(2);
    Operation_IFC mod_29_inner = mod_29_bufferize.operation;
    Operation_IFC mod_29 <- mkDebugOperation(mod_29_inner, "mod_29");
    Operation_IFC mod_30_inner <- mkRepeatStatic(8);
    Operation_IFC mod_30 <- mkDebugOperation(mod_30_inner, "mod_30");
    Operation_IFC mod_31_inner <- mkFlatten(1);
    Operation_IFC mod_31 <- mkDebugOperation(mod_31_inner, "mod_31");
    Operation_IFC mod_32_inner <- mkFlatten(0);
    Operation_IFC mod_32 <- mkDebugOperation(mod_32_inner, "mod_32");
    Operation_IFC mod_33_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_33 <- mkDebugOperation(mod_33_inner, "mod_33");
    PMU_IFC mod_34_bufferize <- mkPMU(1);
    Operation_IFC mod_34_inner = mod_34_bufferize.operation;
    Operation_IFC mod_34 <- mkDebugOperation(mod_34_inner, "mod_34");
    Operation_IFC mod_35_inner <- mkRepeatStatic(16);
    Operation_IFC mod_35 <- mkDebugOperation(mod_35_inner, "mod_35");
    PMU_IFC mod_36_bufferize <- mkPMU(2);
    Operation_IFC mod_36_inner = mod_36_bufferize.operation;
    Operation_IFC mod_36 <- mkDebugOperation(mod_36_inner, "mod_36");
    Operation_IFC mod_37_inner <- mkRepeatStatic(8);
    Operation_IFC mod_37 <- mkDebugOperation(mod_37_inner, "mod_37");
    Operation_IFC mod_38_inner <- mkFlatten(1);
    Operation_IFC mod_38 <- mkDebugOperation(mod_38_inner, "mod_38");
    Operation_IFC mod_39_inner <- mkFlatten(0);
    Operation_IFC mod_39 <- mkDebugOperation(mod_39_inner, "mod_39");
    Operation_IFC mod_40_inner <- mkDynamicRandomLoad(Cons(2, Cons(1, Cons(1, Cons(1, Nil)))));
    Operation_IFC mod_40 <- mkDebugOperation(mod_40_inner, "mod_40");
    Operation_IFC mod_41_inner <- mkRepeatStatic(16);
    Operation_IFC mod_41 <- mkDebugOperation(mod_41_inner, "mod_41");
    Operation_IFC mod_42_inner <- mkRepeatStatic(2);
    Operation_IFC mod_42 <- mkDebugOperation(mod_42_inner, "mod_42");
    PMU_IFC mod_43_bufferize <- mkPMU(2);
    Operation_IFC mod_43_inner = mod_43_bufferize.operation;
    Operation_IFC mod_43 <- mkDebugOperation(mod_43_inner, "mod_43");
    rule rule_1;
        ChannelMessage t;
        t <- mod_34.get(1);
        mod_28.put(0, t);
    endrule
    rule rule_2;
        ChannelMessage t;
        t <- mod_43.get(1);
        mod_4.put(1, t);
    endrule
    rule rule_3;
        ChannelMessage t;
        t <- mod_4.get(1);
        mod_5.put(0, t);
    endrule
    rule rule_4;
        ChannelMessage t;
        t <- mod_5.get(1);
        mod_33.put(0, t);
    endrule
    rule rule_5;
        ChannelMessage t;
        t <- mod_32.get(0);
        mod_31.put(0, t);
    endrule
    rule rule_6;
        ChannelMessage t;
        t <- mod_29.get(1);
        mod_28.put(1, t);
    endrule
    rule rule_7;
        ChannelMessage t;
        t <- mod_14.get(0);
        mod_15.put(0, t);
    endrule
    rule rule_8;
        ChannelMessage t;
        t <- mod_37.get(0);
        mod_36.put(1, t);
    endrule
    rule rule_9;
        ChannelMessage t;
        t <- mod_8.get(0);
        mod_41.put(0, t);
    endrule
    rule rule_10;
        ChannelMessage t;
        t <- mod_12.get(1);
        mod_13.put(0, t);
    endrule
    rule rule_11;
        ChannelMessage t;
        t <- mod_18.get(0);
        mod_18.put(1, t);
    endrule
    rule rule_12;
        ChannelMessage t;
        t <- mod_10.get(0);
        mod_11.put(0, t);
    endrule
    rule rule_13;
        ChannelMessage t;
        t <- mod_9.get(0);
        mod_10.put(0, t);
    endrule
    rule rule_14;
        ChannelMessage t;
        t <- mod_20.get(1);
        mod_13.put(1, t);
    endrule
    rule rule_15;
        ChannelMessage t;
        t <- mod_11.get(0);
        mod_12.put(0, t);
    endrule
    rule rule_16;
        ChannelMessage t;
        t <- mod_28.get(0);
        mod_27.put(0, t);
    endrule
    rule rule_17;
        ChannelMessage t;
        t <- mod_16.get(0);
        mod_18.put(0, t);
    endrule
    rule rule_18;
        ChannelMessage t;
        t <- mod_20.get(0);
        mod_21.put(0, t);
    endrule
    rule rule_19;
        ChannelMessage t;
        t <- mod_2.get(0);
        mod_3.put(0, t);
    endrule
    rule rule_20;
        ChannelMessage t;
        t <- mod_19.get(1);
        mod_15.put(1, t);
    endrule
    rule rule_21;
        ChannelMessage t;
        t <- mod_38.get(0);
        mod_36.put(0, t);
    endrule
    rule rule_22;
        ChannelMessage t;
        t <- mod_7.get(0);
        mod_34.put(0, t);
    endrule
    rule rule_23;
        ChannelMessage t;
        t <- mod_21.get(0);
        mod_20.put(1, t);
    endrule
    rule rule_24;
        ChannelMessage t;
        t <- mod_34.get(0);
        mod_35.put(0, t);
    endrule
    rule rule_25;
        ChannelMessage t;
        t <- mod_36.get(0);
        mod_37.put(0, t);
    endrule
    rule rule_26;
        ChannelMessage t;
        t <- mod_42.get(0);
        mod_6.put(1, t);
    endrule
    rule rule_27;
        ChannelMessage t;
        t <- mod_30.get(0);
        mod_29.put(1, t);
    endrule
    rule rule_28;
        ChannelMessage t;
        t <- mod_23.get(0);
        mod_22.put(0, t);
    endrule
    rule rule_29;
        ChannelMessage t;
        t <- mod_27.get(0);
        mod_26.put(0, t);
    endrule
    rule rule_30;
        ChannelMessage t;
        t <- mod_36.get(1);
        mod_9.put(1, t);
    endrule
    rule rule_31;
        ChannelMessage t;
        t <- mod_15.get(0);
        mod_19.put(0, t);
    endrule
    rule rule_32;
        ChannelMessage t;
        t <- mod_33.get(0);
        mod_32.put(0, t);
    endrule
    rule rule_33;
        ChannelMessage t;
        t <- mod_35.get(0);
        mod_34.put(1, t);
    endrule
    rule rule_34;
        ChannelMessage t;
        t <- mod_6.get(0);
        mod_42.put(0, t);
    endrule
    rule rule_35;
        ChannelMessage t;
        t <- mod_4.get(0);
        mod_43.put(0, t);
    endrule
    rule rule_36;
        ChannelMessage t;
        t <- mod_25.get(0);
        mod_12.put(1, t);
    endrule
    rule rule_37;
        ChannelMessage t;
        t <- mod_16.get(1);
        mod_17.put(1, t);
    endrule
    rule rule_38;
        ChannelMessage t;
        t <- mod_8.get(1);
        mod_9.put(0, t);
    endrule
    rule rule_39;
        ChannelMessage t;
        t <- mod_15.get(1);
        mod_16.put(0, t);
    endrule
    rule rule_40;
        ChannelMessage t;
        t <- mod_5.get(0);
        mod_24.put(0, t);
    endrule
    rule rule_41;
        ChannelMessage t;
        t <- mod_18.get(1);
        mod_16.put(1, t);
    endrule
    rule rule_42;
        ChannelMessage t;
        t <- mod_1.get(0);
        mod_2.put(0, t);
    endrule
    rule rule_43;
        ChannelMessage t;
        t <- mod_12.get(0);
        mod_25.put(0, t);
    endrule
    rule rule_44;
        ChannelMessage t;
        t <- mod_5.get(3);
        mod_6.put(0, t);
    endrule
    rule rule_45;
        ChannelMessage t;
        t <- mod_5.get(2);
        mod_40.put(0, t);
    endrule
    rule rule_46;
        ChannelMessage t;
        t <- mod_19.get(0);
        mod_19.put(1, t);
    endrule
    rule rule_47;
        ChannelMessage t;
        t <- mod_26.get(0);
        mod_11.put(1, t);
    endrule
    rule rule_48;
        ChannelMessage t;
        t <- mod_29.get(0);
        mod_30.put(0, t);
    endrule
    rule rule_49;
        ChannelMessage t;
        t <- mod_31.get(0);
        mod_29.put(0, t);
    endrule
    rule rule_50;
        ChannelMessage t;
        t <- mod_40.get(0);
        mod_39.put(0, t);
    endrule
    rule rule_51;
        ChannelMessage t;
        t <- mod_6.get(1);
        mod_7.put(0, t);
    endrule
    rule rule_52;
        ChannelMessage t;
        t <- mod_7.get(1);
        mod_8.put(0, t);
    endrule
    rule rule_53;
        ChannelMessage t;
        t <- mod_41.get(0);
        mod_8.put(1, t);
    endrule
    rule rule_54;
        ChannelMessage t;
        t <- mod_13.get(0);
        mod_14.put(0, t);
    endrule
    rule rule_55;
        ChannelMessage t;
        t <- mod_24.get(0);
        mod_23.put(0, t);
    endrule
    rule rule_56;
        ChannelMessage t;
        t <- mod_39.get(0);
        mod_38.put(0, t);
    endrule
    rule rule_57;
        ChannelMessage t;
        t <- mod_43.get(0);
        mod_43.put(1, t);
    endrule
    rule rule_58;
        ChannelMessage t;
        t <- mod_3.get(0);
        mod_4.put(0, t);
    endrule
    rule rule_59;
        ChannelMessage t;
        t <- mod_22.get(0);
        mod_20.put(0, t);
    endrule
    method Action put(Int#(32) i, ChannelMessage t);
        if (i == 0) begin
            mod_1.put(0, t);
        end
        if (i == 1) begin
            mod_17.put(0, t);
        end

    endmethod
    method ActionValue#(ChannelMessage) get(Int#(32) i);
        ChannelMessage t = unpack(0);
        if (i == 0) begin
            t <- mod_17.get(0);
        end

        return t;
    endmethod
endmodule

module mkStep(Empty);
    Operation_IFC mod_0_inner <- mkHypernode;
    Operation_IFC mod_0 <- mkDebugOperation(mod_0_inner, "mod_0");
    Operation_IFC mod_44_inner <- mkHypernode;
    Operation_IFC mod_44 <- mkDebugOperation(mod_44_inner, "mod_44");
    Operation_IFC mod_88_inner <- mkHypernode;
    Operation_IFC mod_88 <- mkDebugOperation(mod_88_inner, "mod_88");
    Operation_IFC mod_132_inner <- mkHypernode;
    Operation_IFC mod_132 <- mkDebugOperation(mod_132_inner, "mod_132");
    Operation_IFC mod_176_inner <- mkHypernode;
    Operation_IFC mod_176 <- mkDebugOperation(mod_176_inner, "mod_176");
    Operation_IFC mod_220_inner <- mkHypernode;
    Operation_IFC mod_220 <- mkDebugOperation(mod_220_inner, "mod_220");
    Operation_IFC mod_264_inner <- mkHypernode;
    Operation_IFC mod_264 <- mkDebugOperation(mod_264_inner, "mod_264");
    Operation_IFC mod_308_inner <- mkHypernode;
    Operation_IFC mod_308 <- mkDebugOperation(mod_308_inner, "mod_308");
    Operation_IFC mod_352_inner <- mkHypernode;
    Operation_IFC mod_352 <- mkDebugOperation(mod_352_inner, "mod_352");
    Operation_IFC mod_396_inner <- mkHypernode;
    Operation_IFC mod_396 <- mkDebugOperation(mod_396_inner, "mod_396");
    Operation_IFC mod_440_inner <- mkHypernode;
    Operation_IFC mod_440 <- mkDebugOperation(mod_440_inner, "mod_440");
    Operation_IFC mod_484_inner <- mkHypernode;
    Operation_IFC mod_484 <- mkDebugOperation(mod_484_inner, "mod_484");
    Operation_IFC mod_528_inner <- mkHypernode;
    Operation_IFC mod_528 <- mkDebugOperation(mod_528_inner, "mod_528");
    Operation_IFC mod_572_inner <- mkHypernode;
    Operation_IFC mod_572 <- mkDebugOperation(mod_572_inner, "mod_572");
    Operation_IFC mod_616_inner <- mkHypernode;
    Operation_IFC mod_616 <- mkDebugOperation(mod_616_inner, "mod_616");
    Operation_IFC mod_660_inner <- mkHypernode;
    Operation_IFC mod_660 <- mkDebugOperation(mod_660_inner, "mod_660");
    Operation_IFC mod_704_inner <- mkHypernode;
    Operation_IFC mod_704 <- mkDebugOperation(mod_704_inner, "mod_704");
    Operation_IFC mod_748_inner <- mkHypernode;
    Operation_IFC mod_748 <- mkDebugOperation(mod_748_inner, "mod_748");
    Operation_IFC mod_792_inner <- mkHypernode;
    Operation_IFC mod_792 <- mkDebugOperation(mod_792_inner, "mod_792");
    Operation_IFC mod_836_inner <- mkHypernode;
    Operation_IFC mod_836 <- mkDebugOperation(mod_836_inner, "mod_836");
    Operation_IFC mod_880_inner <- mkHypernode;
    Operation_IFC mod_880 <- mkDebugOperation(mod_880_inner, "mod_880");
    Operation_IFC mod_924_inner <- mkHypernode;
    Operation_IFC mod_924 <- mkDebugOperation(mod_924_inner, "mod_924");
    Operation_IFC mod_968_inner <- mkHypernode;
    Operation_IFC mod_968 <- mkDebugOperation(mod_968_inner, "mod_968");
    Operation_IFC mod_1012_inner <- mkHypernode;
    Operation_IFC mod_1012 <- mkDebugOperation(mod_1012_inner, "mod_1012");
    Operation_IFC mod_1056_inner <- mkHypernode;
    Operation_IFC mod_1056 <- mkDebugOperation(mod_1056_inner, "mod_1056");
    Operation_IFC mod_1100_inner <- mkHypernode;
    Operation_IFC mod_1100 <- mkDebugOperation(mod_1100_inner, "mod_1100");
    Operation_IFC mod_1144_inner <- mkHypernode;
    Operation_IFC mod_1144 <- mkDebugOperation(mod_1144_inner, "mod_1144");
    Operation_IFC mod_1188_inner <- mkHypernode;
    Operation_IFC mod_1188 <- mkDebugOperation(mod_1188_inner, "mod_1188");
    Operation_IFC mod_1232_inner <- mkHypernode;
    Operation_IFC mod_1232 <- mkDebugOperation(mod_1232_inner, "mod_1232");
    Operation_IFC mod_1276_inner <- mkHypernode;
    Operation_IFC mod_1276 <- mkDebugOperation(mod_1276_inner, "mod_1276");
    Operation_IFC mod_1320_inner <- mkHypernode;
    Operation_IFC mod_1320 <- mkDebugOperation(mod_1320_inner, "mod_1320");
    Operation_IFC mod_1364_inner <- mkHypernode;
    Operation_IFC mod_1364 <- mkDebugOperation(mod_1364_inner, "mod_1364");
    Operation_IFC mod_1408_inner <- mkHypernode;
    Operation_IFC mod_1408 <- mkDebugOperation(mod_1408_inner, "mod_1408");
    Operation_IFC mod_1452_inner <- mkHypernode;
    Operation_IFC mod_1452 <- mkDebugOperation(mod_1452_inner, "mod_1452");
    Operation_IFC mod_1496_inner <- mkHypernode;
    Operation_IFC mod_1496 <- mkDebugOperation(mod_1496_inner, "mod_1496");
    Operation_IFC mod_1540_inner <- mkHypernode;
    Operation_IFC mod_1540 <- mkDebugOperation(mod_1540_inner, "mod_1540");
    Operation_IFC mod_1584_inner <- mkHypernode;
    Operation_IFC mod_1584 <- mkDebugOperation(mod_1584_inner, "mod_1584");
    Operation_IFC mod_1628_inner <- mkHypernode;
    Operation_IFC mod_1628 <- mkDebugOperation(mod_1628_inner, "mod_1628");
    Operation_IFC mod_1672_inner <- mkHypernode;
    Operation_IFC mod_1672 <- mkDebugOperation(mod_1672_inner, "mod_1672");
    Operation_IFC mod_1716_inner <- mkHypernode;
    Operation_IFC mod_1716 <- mkDebugOperation(mod_1716_inner, "mod_1716");
    Operation_IFC mod_1760_inner <- mkHypernode;
    Operation_IFC mod_1760 <- mkDebugOperation(mod_1760_inner, "mod_1760");
    Operation_IFC mod_1804_inner <- mkHypernode;
    Operation_IFC mod_1804 <- mkDebugOperation(mod_1804_inner, "mod_1804");
    Operation_IFC mod_1848_inner <- mkHypernode;
    Operation_IFC mod_1848 <- mkDebugOperation(mod_1848_inner, "mod_1848");
    Operation_IFC mod_1892_inner <- mkHypernode;
    Operation_IFC mod_1892 <- mkDebugOperation(mod_1892_inner, "mod_1892");
    Operation_IFC mod_1936_inner <- mkHypernode;
    Operation_IFC mod_1936 <- mkDebugOperation(mod_1936_inner, "mod_1936");
    Operation_IFC mod_1980_inner <- mkHypernode;
    Operation_IFC mod_1980 <- mkDebugOperation(mod_1980_inner, "mod_1980");
    Operation_IFC mod_2024_inner <- mkHypernode;
    Operation_IFC mod_2024 <- mkDebugOperation(mod_2024_inner, "mod_2024");
    Operation_IFC mod_2068_inner <- mkHypernode;
    Operation_IFC mod_2068 <- mkDebugOperation(mod_2068_inner, "mod_2068");
    Operation_IFC mod_2112_inner <- mkHypernode;
    Operation_IFC mod_2112 <- mkDebugOperation(mod_2112_inner, "mod_2112");
    Operation_IFC mod_2156_inner <- mkHypernode;
    Operation_IFC mod_2156 <- mkDebugOperation(mod_2156_inner, "mod_2156");
    Operation_IFC mod_2200_inner <- mkHypernode;
    Operation_IFC mod_2200 <- mkDebugOperation(mod_2200_inner, "mod_2200");
    Operation_IFC mod_2244_inner <- mkHypernode;
    Operation_IFC mod_2244 <- mkDebugOperation(mod_2244_inner, "mod_2244");
    Operation_IFC mod_2288_inner <- mkHypernode;
    Operation_IFC mod_2288 <- mkDebugOperation(mod_2288_inner, "mod_2288");
    Operation_IFC mod_2332_inner <- mkHypernode;
    Operation_IFC mod_2332 <- mkDebugOperation(mod_2332_inner, "mod_2332");
    Operation_IFC mod_2376_inner <- mkHypernode;
    Operation_IFC mod_2376 <- mkDebugOperation(mod_2376_inner, "mod_2376");
    Operation_IFC mod_2420_inner <- mkHypernode;
    Operation_IFC mod_2420 <- mkDebugOperation(mod_2420_inner, "mod_2420");
    Operation_IFC mod_2464_inner <- mkHypernode;
    Operation_IFC mod_2464 <- mkDebugOperation(mod_2464_inner, "mod_2464");
    Operation_IFC mod_2508_inner <- mkHypernode;
    Operation_IFC mod_2508 <- mkDebugOperation(mod_2508_inner, "mod_2508");
    Operation_IFC mod_2552_inner <- mkHypernode;
    Operation_IFC mod_2552 <- mkDebugOperation(mod_2552_inner, "mod_2552");
    Operation_IFC mod_2596_inner <- mkHypernode;
    Operation_IFC mod_2596 <- mkDebugOperation(mod_2596_inner, "mod_2596");
    Operation_IFC mod_2640_inner <- mkHypernode;
    Operation_IFC mod_2640 <- mkDebugOperation(mod_2640_inner, "mod_2640");
    Operation_IFC mod_2684_inner <- mkHypernode;
    Operation_IFC mod_2684 <- mkDebugOperation(mod_2684_inner, "mod_2684");
    Operation_IFC mod_2728_inner <- mkHypernode;
    Operation_IFC mod_2728 <- mkDebugOperation(mod_2728_inner, "mod_2728");
    Operation_IFC mod_2772_inner <- mkHypernode;
    Operation_IFC mod_2772 <- mkDebugOperation(mod_2772_inner, "mod_2772");
    Operation_IFC mod_2816_inner <- mkHypernode;
    Operation_IFC mod_2816 <- mkDebugOperation(mod_2816_inner, "mod_2816");
    Operation_IFC mod_2860_inner <- mkHypernode;
    Operation_IFC mod_2860 <- mkDebugOperation(mod_2860_inner, "mod_2860");
    Operation_IFC mod_2904_inner <- mkHypernode;
    Operation_IFC mod_2904 <- mkDebugOperation(mod_2904_inner, "mod_2904");
    Operation_IFC mod_2948_inner <- mkHypernode;
    Operation_IFC mod_2948 <- mkDebugOperation(mod_2948_inner, "mod_2948");
    Operation_IFC mod_2992_inner <- mkHypernode;
    Operation_IFC mod_2992 <- mkDebugOperation(mod_2992_inner, "mod_2992");
    Operation_IFC mod_3036_inner <- mkHypernode;
    Operation_IFC mod_3036 <- mkDebugOperation(mod_3036_inner, "mod_3036");
    Operation_IFC mod_3080_inner <- mkHypernode;
    Operation_IFC mod_3080 <- mkDebugOperation(mod_3080_inner, "mod_3080");
    Operation_IFC mod_3124_inner <- mkHypernode;
    Operation_IFC mod_3124 <- mkDebugOperation(mod_3124_inner, "mod_3124");
    Operation_IFC mod_3168_inner <- mkHypernode;
    Operation_IFC mod_3168 <- mkDebugOperation(mod_3168_inner, "mod_3168");
    Operation_IFC mod_3212_inner <- mkHypernode;
    Operation_IFC mod_3212 <- mkDebugOperation(mod_3212_inner, "mod_3212");
    Operation_IFC mod_3256_inner <- mkHypernode;
    Operation_IFC mod_3256 <- mkDebugOperation(mod_3256_inner, "mod_3256");
    Operation_IFC mod_3300_inner <- mkHypernode;
    Operation_IFC mod_3300 <- mkDebugOperation(mod_3300_inner, "mod_3300");
    Operation_IFC mod_3344_inner <- mkHypernode;
    Operation_IFC mod_3344 <- mkDebugOperation(mod_3344_inner, "mod_3344");
    Operation_IFC mod_3388_inner <- mkHypernode;
    Operation_IFC mod_3388 <- mkDebugOperation(mod_3388_inner, "mod_3388");
    Operation_IFC mod_3432_inner <- mkHypernode;
    Operation_IFC mod_3432 <- mkDebugOperation(mod_3432_inner, "mod_3432");
    Operation_IFC mod_3476_inner <- mkHypernode;
    Operation_IFC mod_3476 <- mkDebugOperation(mod_3476_inner, "mod_3476");
    Operation_IFC mod_3520_inner <- mkHypernode;
    Operation_IFC mod_3520 <- mkDebugOperation(mod_3520_inner, "mod_3520");
    Operation_IFC mod_3564_inner <- mkHypernode;
    Operation_IFC mod_3564 <- mkDebugOperation(mod_3564_inner, "mod_3564");
    Operation_IFC mod_3608_inner <- mkHypernode;
    Operation_IFC mod_3608 <- mkDebugOperation(mod_3608_inner, "mod_3608");
    Operation_IFC mod_3652_inner <- mkHypernode;
    Operation_IFC mod_3652 <- mkDebugOperation(mod_3652_inner, "mod_3652");
    Operation_IFC mod_3696_inner <- mkHypernode;
    Operation_IFC mod_3696 <- mkDebugOperation(mod_3696_inner, "mod_3696");
    Operation_IFC mod_3740_inner <- mkHypernode;
    Operation_IFC mod_3740 <- mkDebugOperation(mod_3740_inner, "mod_3740");
    Operation_IFC mod_3784_inner <- mkHypernode;
    Operation_IFC mod_3784 <- mkDebugOperation(mod_3784_inner, "mod_3784");
    Operation_IFC mod_3828_inner <- mkHypernode;
    Operation_IFC mod_3828 <- mkDebugOperation(mod_3828_inner, "mod_3828");
    Operation_IFC mod_3872_inner <- mkHypernode;
    Operation_IFC mod_3872 <- mkDebugOperation(mod_3872_inner, "mod_3872");
    Operation_IFC mod_3916_inner <- mkHypernode;
    Operation_IFC mod_3916 <- mkDebugOperation(mod_3916_inner, "mod_3916");
    Operation_IFC mod_3960_inner <- mkHypernode;
    Operation_IFC mod_3960 <- mkDebugOperation(mod_3960_inner, "mod_3960");
    Operation_IFC mod_4004_inner <- mkHypernode;
    Operation_IFC mod_4004 <- mkDebugOperation(mod_4004_inner, "mod_4004");
    Operation_IFC mod_4048_inner <- mkHypernode;
    Operation_IFC mod_4048 <- mkDebugOperation(mod_4048_inner, "mod_4048");
    Operation_IFC mod_4092_inner <- mkHypernode;
    Operation_IFC mod_4092 <- mkDebugOperation(mod_4092_inner, "mod_4092");
    Operation_IFC mod_4136_inner <- mkHypernode;
    Operation_IFC mod_4136 <- mkDebugOperation(mod_4136_inner, "mod_4136");
    Operation_IFC mod_4180_inner <- mkHypernode;
    Operation_IFC mod_4180 <- mkDebugOperation(mod_4180_inner, "mod_4180");
    Operation_IFC mod_4224_inner <- mkHypernode;
    Operation_IFC mod_4224 <- mkDebugOperation(mod_4224_inner, "mod_4224");
    Operation_IFC mod_4268_inner <- mkHypernode;
    Operation_IFC mod_4268 <- mkDebugOperation(mod_4268_inner, "mod_4268");
    Operation_IFC mod_4312_inner <- mkHypernode;
    Operation_IFC mod_4312 <- mkDebugOperation(mod_4312_inner, "mod_4312");
    Operation_IFC mod_4356_inner <- mkHypernode;
    Operation_IFC mod_4356 <- mkDebugOperation(mod_4356_inner, "mod_4356");
    Operation_IFC mod_4400_inner <- mkHypernode;
    Operation_IFC mod_4400 <- mkDebugOperation(mod_4400_inner, "mod_4400");
    Operation_IFC mod_4444_inner <- mkHypernode;
    Operation_IFC mod_4444 <- mkDebugOperation(mod_4444_inner, "mod_4444");
    Operation_IFC mod_4488_inner <- mkHypernode;
    Operation_IFC mod_4488 <- mkDebugOperation(mod_4488_inner, "mod_4488");
    Operation_IFC mod_4532_inner <- mkHypernode;
    Operation_IFC mod_4532 <- mkDebugOperation(mod_4532_inner, "mod_4532");
    Operation_IFC mod_4576_inner <- mkHypernode;
    Operation_IFC mod_4576 <- mkDebugOperation(mod_4576_inner, "mod_4576");
    Operation_IFC mod_4620_inner <- mkHypernode;
    Operation_IFC mod_4620 <- mkDebugOperation(mod_4620_inner, "mod_4620");
    Operation_IFC mod_4664_inner <- mkHypernode;
    Operation_IFC mod_4664 <- mkDebugOperation(mod_4664_inner, "mod_4664");
    Operation_IFC mod_4708_inner <- mkHypernode;
    Operation_IFC mod_4708 <- mkDebugOperation(mod_4708_inner, "mod_4708");
    Operation_IFC mod_4752_inner <- mkHypernode;
    Operation_IFC mod_4752 <- mkDebugOperation(mod_4752_inner, "mod_4752");
    Operation_IFC mod_4796_inner <- mkHypernode;
    Operation_IFC mod_4796 <- mkDebugOperation(mod_4796_inner, "mod_4796");
    Operation_IFC mod_4840_inner <- mkHypernode;
    Operation_IFC mod_4840 <- mkDebugOperation(mod_4840_inner, "mod_4840");
    Operation_IFC mod_4884_inner <- mkHypernode;
    Operation_IFC mod_4884 <- mkDebugOperation(mod_4884_inner, "mod_4884");
    Operation_IFC mod_4928_inner <- mkHypernode;
    Operation_IFC mod_4928 <- mkDebugOperation(mod_4928_inner, "mod_4928");
    Operation_IFC mod_4972_inner <- mkHypernode;
    Operation_IFC mod_4972 <- mkDebugOperation(mod_4972_inner, "mod_4972");
    Operation_IFC mod_5016_inner <- mkHypernode;
    Operation_IFC mod_5016 <- mkDebugOperation(mod_5016_inner, "mod_5016");
    Operation_IFC mod_5060_inner <- mkHypernode;
    Operation_IFC mod_5060 <- mkDebugOperation(mod_5060_inner, "mod_5060");
    Operation_IFC mod_5104_inner <- mkHypernode;
    Operation_IFC mod_5104 <- mkDebugOperation(mod_5104_inner, "mod_5104");
    Operation_IFC mod_5148_inner <- mkHypernode;
    Operation_IFC mod_5148 <- mkDebugOperation(mod_5148_inner, "mod_5148");
    Operation_IFC mod_5192_inner <- mkHypernode;
    Operation_IFC mod_5192 <- mkDebugOperation(mod_5192_inner, "mod_5192");
    Operation_IFC mod_5236_inner <- mkHypernode;
    Operation_IFC mod_5236 <- mkDebugOperation(mod_5236_inner, "mod_5236");
    Operation_IFC mod_5280_inner <- mkHypernode;
    Operation_IFC mod_5280 <- mkDebugOperation(mod_5280_inner, "mod_5280");
    Operation_IFC mod_5324_inner <- mkHypernode;
    Operation_IFC mod_5324 <- mkDebugOperation(mod_5324_inner, "mod_5324");
    Operation_IFC mod_5368_inner <- mkHypernode;
    Operation_IFC mod_5368 <- mkDebugOperation(mod_5368_inner, "mod_5368");
    Operation_IFC mod_5412_inner <- mkHypernode;
    Operation_IFC mod_5412 <- mkDebugOperation(mod_5412_inner, "mod_5412");
    Operation_IFC mod_5456_inner <- mkHypernode;
    Operation_IFC mod_5456 <- mkDebugOperation(mod_5456_inner, "mod_5456");
    Operation_IFC mod_5500_inner <- mkHypernode;
    Operation_IFC mod_5500 <- mkDebugOperation(mod_5500_inner, "mod_5500");
    Operation_IFC mod_5544_inner <- mkHypernode;
    Operation_IFC mod_5544 <- mkDebugOperation(mod_5544_inner, "mod_5544");
    Operation_IFC mod_5588_inner <- mkHypernode;
    Operation_IFC mod_5588 <- mkDebugOperation(mod_5588_inner, "mod_5588");
    Operation_IFC mod_5632_inner <- mkRandomOffChipLoad(Cons(64, Cons(1, Cons(1, Cons(1, Cons(1, Cons(1, Nil)))))));
    Operation_IFC mod_5632 <- mkDebugOperation(mod_5632_inner, "mod_5632");
    Partition_IFC#(128) mod_5633_inner <- mkPartition(0, 128);
    Operation_IFC mod_5633 <- mkDebugOperation(mod_5633_inner.op, "mod_5633");
    Partition_IFC#(128) mod_5634_inner <- mkPartition(0, 128);
    Operation_IFC mod_5634 <- mkDebugOperation(mod_5634_inner.op, "mod_5634");
    Reassemble_IFC#(128) mod_5635_inner <- mkReassemble(128);
    Operation_IFC mod_5635 <- mkDebugOperation(mod_5635_inner.op, "mod_5635");
    Operation_IFC mod_5636_inner <- mkFlatten(1);
    Operation_IFC mod_5636 <- mkDebugOperation(mod_5636_inner, "mod_5636");
    Operation_IFC mod_5637_inner <- mkReshape(2, 1);
    Operation_IFC mod_5637 <- mkDebugOperation(mod_5637_inner, "mod_5637");
    PMU_IFC mod_5638_bufferize <- mkPMU(2);
    Operation_IFC mod_5638_inner = mod_5638_bufferize.operation;
    Operation_IFC mod_5638 <- mkDebugOperation(mod_5638_inner, "mod_5638");
    Operation_IFC mod_5639_inner <- mkRepeatStatic(1);
    Operation_IFC mod_5639 <- mkDebugOperation(mod_5639_inner, "mod_5639");
    Operation_IFC mod_5640_inner <- mkRandomSelectGen(128);
    Operation_IFC mod_5640 <- mkDebugOperation(mod_5640_inner, "mod_5640");
    Operation_IFC mod_5641_inner <- mkPrinter("mod_5641");
    Operation_IFC mod_5641 <- mkDebugOperation(mod_5641_inner, "mod_5641");
    Operation_IFC mod_5642_inner <- mkFlatten(0);
    Operation_IFC mod_5642 <- mkDebugOperation(mod_5642_inner, "mod_5642");
    Operation_IFC mod_5643_inner <- mkRepeatStatic(1);
    Operation_IFC mod_5643 <- mkDebugOperation(mod_5643_inner, "mod_5643");
    Operation_IFC mod_5644_inner <- mkRandomOffChipLoad(Cons(64, Cons(8, Cons(1, Cons(1, Cons(1, Cons(1, Nil)))))));
    Operation_IFC mod_5644 <- mkDebugOperation(mod_5644_inner, "mod_5644");
    Operation_IFC mod_5645_inner <- mkAccumBigTile(add_tile, 3);
    Operation_IFC mod_5645 <- mkDebugOperation(mod_5645_inner, "mod_5645");
    Operation_IFC mod_5646_inner <- mkRepeatStatic(1);
    Operation_IFC mod_5646 <- mkDebugOperation(mod_5646_inner, "mod_5646");
    Operation_IFC mod_5647_inner <- mkRandomSelectGen(128);
    Operation_IFC mod_5647 <- mkDebugOperation(mod_5647_inner, "mod_5647");
    Operation_IFC mod_5648_inner <- mkRandomSelectGen(128);
    Operation_IFC mod_5648 <- mkDebugOperation(mod_5648_inner, "mod_5648");
    (* descending_urgency = "rule_1, rule_2, rule_3, rule_4, rule_5, rule_6, rule_7, rule_8, rule_9, rule_10, rule_11, rule_12, rule_13, rule_14, rule_15, rule_16, rule_17, rule_18, rule_19, rule_20, rule_21, rule_22, rule_23, rule_24, rule_25, rule_26, rule_27, rule_28, rule_29, rule_30, rule_31, rule_32, rule_33, rule_34, rule_35, rule_36, rule_37, rule_38, rule_39, rule_40, rule_41, rule_42, rule_43, rule_44, rule_45, rule_46, rule_47, rule_48, rule_49, rule_50, rule_51, rule_52, rule_53, rule_54, rule_55, rule_56, rule_57, rule_58, rule_59, rule_60, rule_61, rule_62, rule_63, rule_64, rule_65, rule_66, rule_67, rule_68, rule_69, rule_70, rule_71, rule_72, rule_73, rule_74, rule_75, rule_76, rule_77, rule_78, rule_79, rule_80, rule_81, rule_82, rule_83, rule_84, rule_85, rule_86, rule_87, rule_88, rule_89, rule_90, rule_91, rule_92, rule_93, rule_94, rule_95, rule_96, rule_97, rule_98, rule_99, rule_100, rule_101, rule_102, rule_103, rule_104, rule_105, rule_106, rule_107, rule_108, rule_109, rule_110, rule_111, rule_112, rule_113, rule_114, rule_115, rule_116, rule_117, rule_118, rule_119, rule_120, rule_121, rule_122, rule_123, rule_124, rule_125, rule_126, rule_127, rule_128, rule_129, rule_130, rule_131, rule_132, rule_133, rule_134, rule_135, rule_136, rule_137, rule_138, rule_139, rule_140, rule_141, rule_142, rule_143, rule_144, rule_145, rule_146, rule_147, rule_148, rule_149, rule_150, rule_151, rule_152, rule_153, rule_154, rule_155, rule_156, rule_157, rule_158, rule_159, rule_160, rule_161, rule_162, rule_163, rule_164, rule_165, rule_166, rule_167, rule_168, rule_169, rule_170, rule_171, rule_172, rule_173, rule_174, rule_175, rule_176, rule_177, rule_178, rule_179, rule_180, rule_181, rule_182, rule_183, rule_184, rule_185, rule_186, rule_187, rule_188, rule_189, rule_190, rule_191, rule_192, rule_193, rule_194, rule_195, rule_196, rule_197, rule_198, rule_199, rule_200, rule_201, rule_202, rule_203, rule_204, rule_205, rule_206, rule_207, rule_208, rule_209, rule_210, rule_211, rule_212, rule_213, rule_214, rule_215, rule_216, rule_217, rule_218, rule_219, rule_220, rule_221, rule_222, rule_223, rule_224, rule_225, rule_226, rule_227, rule_228, rule_229, rule_230, rule_231, rule_232, rule_233, rule_234, rule_235, rule_236, rule_237, rule_238, rule_239, rule_240, rule_241, rule_242, rule_243, rule_244, rule_245, rule_246, rule_247, rule_248, rule_249, rule_250, rule_251, rule_252, rule_253, rule_254, rule_255, rule_256, rule_257, rule_258, rule_259, rule_260, rule_261, rule_262, rule_263, rule_264, rule_265, rule_266, rule_267, rule_268, rule_269, rule_270, rule_271, rule_272, rule_273, rule_274, rule_275, rule_276, rule_277, rule_278, rule_279, rule_280, rule_281, rule_282, rule_283, rule_284, rule_285, rule_286, rule_287, rule_288, rule_289, rule_290, rule_291, rule_292, rule_293, rule_294, rule_295, rule_296, rule_297, rule_298, rule_299, rule_300, rule_301, rule_302, rule_303, rule_304, rule_305, rule_306, rule_307, rule_308, rule_309, rule_310, rule_311, rule_312, rule_313, rule_314, rule_315, rule_316, rule_317, rule_318, rule_319, rule_320, rule_321, rule_322, rule_323, rule_324, rule_325, rule_326, rule_327, rule_328, rule_329, rule_330, rule_331, rule_332, rule_333, rule_334, rule_335, rule_336, rule_337, rule_338, rule_339, rule_340, rule_341, rule_342, rule_343, rule_344, rule_345, rule_346, rule_347, rule_348, rule_349, rule_350, rule_351, rule_352, rule_353, rule_354, rule_355, rule_356, rule_357, rule_358, rule_359, rule_360, rule_361, rule_362, rule_363, rule_364, rule_365, rule_366, rule_367, rule_368, rule_369, rule_370, rule_371, rule_372, rule_373, rule_374, rule_375, rule_376, rule_377, rule_378, rule_379, rule_380, rule_381, rule_382, rule_383, rule_384, rule_385, rule_386, rule_387, rule_388, rule_389, rule_390, rule_391, rule_392, rule_393, rule_394, rule_395, rule_396, rule_397, rule_398, rule_399, rule_400" *)
    rule rule_1;
        ChannelMessage t;
        t <- mod_5633.get(20);
        mod_880.put(1, t);
    endrule
    rule rule_2;
        ChannelMessage t;
        t <- mod_1320.get(0);
        mod_5635.put(97, t);
    endrule
    rule rule_3;
        ChannelMessage t;
        t <- mod_5633.get(122);
        mod_5368.put(1, t);
    endrule
    rule rule_4;
        ChannelMessage t;
        t <- mod_5634.get(64);
        mod_2816.put(0, t);
    endrule
    rule rule_5;
        ChannelMessage t;
        t <- mod_5633.get(55);
        mod_2420.put(1, t);
    endrule
    rule rule_6;
        ChannelMessage t;
        t <- mod_5634.get(18);
        mod_792.put(0, t);
    endrule
    rule rule_7;
        ChannelMessage t;
        t <- mod_1628.get(0);
        mod_5635.put(90, t);
    endrule
    rule rule_8;
        ChannelMessage t;
        t <- mod_836.get(0);
        mod_5635.put(108, t);
    endrule
    rule rule_9;
        ChannelMessage t;
        t <- mod_3036.get(0);
        mod_5635.put(58, t);
    endrule
    rule rule_10;
        ChannelMessage t;
        t <- mod_4400.get(0);
        mod_5635.put(27, t);
    endrule
    rule rule_11;
        ChannelMessage t;
        t <- mod_5633.get(53);
        mod_2332.put(1, t);
    endrule
    rule rule_12;
        ChannelMessage t;
        t <- mod_5633.get(82);
        mod_3608.put(1, t);
    endrule
    rule rule_13;
        ChannelMessage t;
        t <- mod_5633.get(21);
        mod_924.put(1, t);
    endrule
    rule rule_14;
        ChannelMessage t;
        t <- mod_5633.get(0);
        mod_0.put(1, t);
    endrule
    rule rule_15;
        ChannelMessage t;
        t <- mod_5633.get(50);
        mod_2200.put(1, t);
    endrule
    rule rule_16;
        ChannelMessage t;
        t <- mod_5634.get(7);
        mod_308.put(0, t);
    endrule
    rule rule_17;
        ChannelMessage t;
        t <- mod_5634.get(62);
        mod_2728.put(0, t);
    endrule
    rule rule_18;
        ChannelMessage t;
        t <- mod_2640.get(0);
        mod_5635.put(67, t);
    endrule
    rule rule_19;
        ChannelMessage t;
        t <- mod_2200.get(0);
        mod_5635.put(77, t);
    endrule
    rule rule_20;
        ChannelMessage t;
        t <- mod_5633.get(19);
        mod_836.put(1, t);
    endrule
    rule rule_21;
        ChannelMessage t;
        t <- mod_5633.get(37);
        mod_1628.put(1, t);
    endrule
    rule rule_22;
        ChannelMessage t;
        t <- mod_5634.get(74);
        mod_3256.put(0, t);
    endrule
    rule rule_23;
        ChannelMessage t;
        t <- mod_5634.get(127);
        mod_5588.put(0, t);
    endrule
    rule rule_24;
        ChannelMessage t;
        t <- mod_3828.get(0);
        mod_5635.put(40, t);
    endrule
    rule rule_25;
        ChannelMessage t;
        t <- mod_5634.get(16);
        mod_704.put(0, t);
    endrule
    rule rule_26;
        ChannelMessage t;
        t <- mod_5634.get(25);
        mod_1100.put(0, t);
    endrule
    rule rule_27;
        ChannelMessage t;
        t <- mod_5633.get(13);
        mod_572.put(1, t);
    endrule
    rule rule_28;
        ChannelMessage t;
        t <- mod_5633.get(58);
        mod_2552.put(1, t);
    endrule
    rule rule_29;
        ChannelMessage t;
        t <- mod_5633.get(112);
        mod_4928.put(1, t);
    endrule
    rule rule_30;
        ChannelMessage t;
        t <- mod_2992.get(0);
        mod_5635.put(59, t);
    endrule
    rule rule_31;
        ChannelMessage t;
        t <- mod_5634.get(109);
        mod_4796.put(0, t);
    endrule
    rule rule_32;
        ChannelMessage t;
        t <- mod_4356.get(0);
        mod_5635.put(28, t);
    endrule
    rule rule_33;
        ChannelMessage t;
        t <- mod_5633.get(111);
        mod_4884.put(1, t);
    endrule
    rule rule_34;
        ChannelMessage t;
        t <- mod_5634.get(117);
        mod_5148.put(0, t);
    endrule
    rule rule_35;
        ChannelMessage t;
        t <- mod_5634.get(10);
        mod_440.put(0, t);
    endrule
    rule rule_36;
        ChannelMessage t;
        t <- mod_5633.get(92);
        mod_4048.put(1, t);
    endrule
    rule rule_37;
        ChannelMessage t;
        t <- mod_5633.get(25);
        mod_1100.put(1, t);
    endrule
    rule rule_38;
        ChannelMessage t;
        t <- mod_5633.get(102);
        mod_4488.put(1, t);
    endrule
    rule rule_39;
        ChannelMessage t;
        t <- mod_5633.get(73);
        mod_3212.put(1, t);
    endrule
    rule rule_40;
        ChannelMessage t;
        t <- mod_5634.get(93);
        mod_4092.put(0, t);
    endrule
    rule rule_41;
        ChannelMessage t;
        t <- mod_3916.get(0);
        mod_5635.put(38, t);
    endrule
    rule rule_42;
        ChannelMessage t;
        t <- mod_5633.get(70);
        mod_3080.put(1, t);
    endrule
    rule rule_43;
        ChannelMessage t;
        t <- mod_5633.get(86);
        mod_3784.put(1, t);
    endrule
    rule rule_44;
        ChannelMessage t;
        t <- mod_5634.get(106);
        mod_4664.put(0, t);
    endrule
    rule rule_45;
        ChannelMessage t;
        t <- mod_5633.get(63);
        mod_2772.put(1, t);
    endrule
    rule rule_46;
        ChannelMessage t;
        t <- mod_5634.get(94);
        mod_4136.put(0, t);
    endrule
    rule rule_47;
        ChannelMessage t;
        t <- mod_2420.get(0);
        mod_5635.put(72, t);
    endrule
    rule rule_48;
        ChannelMessage t;
        t <- mod_5633.get(31);
        mod_1364.put(1, t);
    endrule
    rule rule_49;
        ChannelMessage t;
        t <- mod_5634.get(68);
        mod_2992.put(0, t);
    endrule
    rule rule_50;
        ChannelMessage t;
        t <- mod_3696.get(0);
        mod_5635.put(43, t);
    endrule
    rule rule_51;
        ChannelMessage t;
        t <- mod_5634.get(49);
        mod_2156.put(0, t);
    endrule
    rule rule_52;
        ChannelMessage t;
        t <- mod_5642.get(0);
        mod_5636.put(0, t);
    endrule
    rule rule_53;
        ChannelMessage t;
        t <- mod_5633.get(72);
        mod_3168.put(1, t);
    endrule
    rule rule_54;
        ChannelMessage t;
        t <- mod_2904.get(0);
        mod_5635.put(61, t);
    endrule
    rule rule_55;
        ChannelMessage t;
        t <- mod_4312.get(0);
        mod_5635.put(29, t);
    endrule
    rule rule_56;
        ChannelMessage t;
        t <- mod_5633.get(12);
        mod_528.put(1, t);
    endrule
    rule rule_57;
        ChannelMessage t;
        t <- mod_5633.get(28);
        mod_1232.put(1, t);
    endrule
    rule rule_58;
        ChannelMessage t;
        t <- mod_5633.get(80);
        mod_3520.put(1, t);
    endrule
    rule rule_59;
        ChannelMessage t;
        t <- mod_5634.get(30);
        mod_1320.put(0, t);
    endrule
    rule rule_60;
        ChannelMessage t;
        t <- mod_1804.get(0);
        mod_5635.put(86, t);
    endrule
    rule rule_61;
        ChannelMessage t;
        t <- mod_5634.get(0);
        mod_0.put(0, t);
    endrule
    rule rule_62;
        ChannelMessage t;
        t <- mod_5634.get(47);
        mod_2068.put(0, t);
    endrule
    rule rule_63;
        ChannelMessage t;
        t <- mod_5634.get(54);
        mod_2376.put(0, t);
    endrule
    rule rule_64;
        ChannelMessage t;
        t <- mod_5634.get(107);
        mod_4708.put(0, t);
    endrule
    rule rule_65;
        ChannelMessage t;
        t <- mod_5645.get(1);
        mod_5637.put(0, t);
    endrule
    rule rule_66;
        ChannelMessage t;
        t <- mod_5634.get(66);
        mod_2904.put(0, t);
    endrule
    rule rule_67;
        ChannelMessage t;
        t <- mod_5634.get(115);
        mod_5060.put(0, t);
    endrule
    rule rule_68;
        ChannelMessage t;
        t <- mod_484.get(0);
        mod_5635.put(116, t);
    endrule
    rule rule_69;
        ChannelMessage t;
        t <- mod_1056.get(0);
        mod_5635.put(103, t);
    endrule
    rule rule_70;
        ChannelMessage t;
        t <- mod_2112.get(0);
        mod_5635.put(79, t);
    endrule
    rule rule_71;
        ChannelMessage t;
        t <- mod_5633.get(49);
        mod_2156.put(1, t);
    endrule
    rule rule_72;
        ChannelMessage t;
        t <- mod_2024.get(0);
        mod_5635.put(81, t);
    endrule
    rule rule_73;
        ChannelMessage t;
        t <- mod_5633.get(95);
        mod_4180.put(1, t);
    endrule
    rule rule_74;
        ChannelMessage t;
        t <- mod_4048.get(0);
        mod_5635.put(35, t);
    endrule
    rule rule_75;
        ChannelMessage t;
        t <- mod_5633.get(68);
        mod_2992.put(1, t);
    endrule
    rule rule_76;
        ChannelMessage t;
        t <- mod_5544.get(0);
        mod_5635.put(1, t);
    endrule
    rule rule_77;
        ChannelMessage t;
        t <- mod_5633.get(71);
        mod_3124.put(1, t);
    endrule
    rule rule_78;
        ChannelMessage t;
        t <- mod_5633.get(118);
        mod_5192.put(1, t);
    endrule
    rule rule_79;
        ChannelMessage t;
        t <- mod_3608.get(0);
        mod_5635.put(45, t);
    endrule
    rule rule_80;
        ChannelMessage t;
        t <- mod_528.get(0);
        mod_5635.put(115, t);
    endrule
    rule rule_81;
        ChannelMessage t;
        t <- mod_2288.get(0);
        mod_5635.put(75, t);
    endrule
    rule rule_82;
        ChannelMessage t;
        t <- mod_2332.get(0);
        mod_5635.put(74, t);
    endrule
    rule rule_83;
        ChannelMessage t;
        t <- mod_5634.get(72);
        mod_3168.put(0, t);
    endrule
    rule rule_84;
        ChannelMessage t;
        t <- mod_5633.get(64);
        mod_2816.put(1, t);
    endrule
    rule rule_85;
        ChannelMessage t;
        t <- mod_5634.get(114);
        mod_5016.put(0, t);
    endrule
    rule rule_86;
        ChannelMessage t;
        t <- mod_5633.get(15);
        mod_660.put(1, t);
    endrule
    rule rule_87;
        ChannelMessage t;
        t <- mod_5634.get(31);
        mod_1364.put(0, t);
    endrule
    rule rule_88;
        ChannelMessage t;
        t <- mod_5633.get(127);
        mod_5588.put(1, t);
    endrule
    rule rule_89;
        ChannelMessage t;
        t <- mod_968.get(0);
        mod_5635.put(105, t);
    endrule
    rule rule_90;
        ChannelMessage t;
        t <- mod_4796.get(0);
        mod_5635.put(18, t);
    endrule
    rule rule_91;
        ChannelMessage t;
        t <- mod_2596.get(0);
        mod_5635.put(68, t);
    endrule
    rule rule_92;
        ChannelMessage t;
        t <- mod_5633.get(105);
        mod_4620.put(1, t);
    endrule
    rule rule_93;
        ChannelMessage t;
        t <- mod_3256.get(0);
        mod_5635.put(53, t);
    endrule
    rule rule_94;
        ChannelMessage t;
        t <- mod_5633.get(113);
        mod_4972.put(1, t);
    endrule
    rule rule_95;
        ChannelMessage t;
        t <- mod_5633.get(103);
        mod_4532.put(1, t);
    endrule
    rule rule_96;
        ChannelMessage t;
        t <- mod_5634.get(85);
        mod_3740.put(0, t);
    endrule
    rule rule_97;
        ChannelMessage t;
        t <- mod_176.get(0);
        mod_5635.put(123, t);
    endrule
    rule rule_98;
        ChannelMessage t;
        t <- mod_3740.get(0);
        mod_5635.put(42, t);
    endrule
    rule rule_99;
        ChannelMessage t;
        t <- mod_308.get(0);
        mod_5635.put(120, t);
    endrule
    rule rule_100;
        ChannelMessage t;
        t <- mod_5236.get(0);
        mod_5635.put(8, t);
    endrule
    rule rule_101;
        ChannelMessage t;
        t <- mod_5633.get(62);
        mod_2728.put(1, t);
    endrule
    rule rule_102;
        ChannelMessage t;
        t <- mod_264.get(0);
        mod_5635.put(121, t);
    endrule
    rule rule_103;
        ChannelMessage t;
        t <- mod_5634.get(28);
        mod_1232.put(0, t);
    endrule
    rule rule_104;
        ChannelMessage t;
        t <- mod_5633.get(7);
        mod_308.put(1, t);
    endrule
    rule rule_105;
        ChannelMessage t;
        t <- mod_5634.get(60);
        mod_2640.put(0, t);
    endrule
    rule rule_106;
        ChannelMessage t;
        t <- mod_5633.get(96);
        mod_4224.put(1, t);
    endrule
    rule rule_107;
        ChannelMessage t;
        t <- mod_3564.get(0);
        mod_5635.put(46, t);
    endrule
    rule rule_108;
        ChannelMessage t;
        t <- mod_5634.get(103);
        mod_4532.put(0, t);
    endrule
    rule rule_109;
        ChannelMessage t;
        t <- mod_5633.get(36);
        mod_1584.put(1, t);
    endrule
    rule rule_110;
        ChannelMessage t;
        t <- mod_5637.get(0);
        mod_5641.put(0, t);
    endrule
    rule rule_111;
        ChannelMessage t;
        t <- mod_5633.get(110);
        mod_4840.put(1, t);
    endrule
    rule rule_112;
        ChannelMessage t;
        t <- mod_5633.get(48);
        mod_2112.put(1, t);
    endrule
    rule rule_113;
        ChannelMessage t;
        t <- mod_5633.get(115);
        mod_5060.put(1, t);
    endrule
    rule rule_114;
        ChannelMessage t;
        t <- mod_5638.get(1);
        mod_5645.put(1, t);
    endrule
    rule rule_115;
        ChannelMessage t;
        t <- mod_4532.get(0);
        mod_5635.put(24, t);
    endrule
    rule rule_116;
        ChannelMessage t;
        t <- mod_5633.get(78);
        mod_3432.put(1, t);
    endrule
    rule rule_117;
        ChannelMessage t;
        t <- mod_2376.get(0);
        mod_5635.put(73, t);
    endrule
    rule rule_118;
        ChannelMessage t;
        t <- mod_1188.get(0);
        mod_5635.put(100, t);
    endrule
    rule rule_119;
        ChannelMessage t;
        t <- mod_5633.get(75);
        mod_3300.put(1, t);
    endrule
    rule rule_120;
        ChannelMessage t;
        t <- mod_3432.get(0);
        mod_5635.put(49, t);
    endrule
    rule rule_121;
        ChannelMessage t;
        t <- mod_5633.get(51);
        mod_2244.put(1, t);
    endrule
    rule rule_122;
        ChannelMessage t;
        t <- mod_5634.get(22);
        mod_968.put(0, t);
    endrule
    rule rule_123;
        ChannelMessage t;
        t <- mod_2156.get(0);
        mod_5635.put(78, t);
    endrule
    rule rule_124;
        ChannelMessage t;
        t <- mod_5632.get(0);
        mod_5642.put(0, t);
    endrule
    rule rule_125;
        ChannelMessage t;
        t <- mod_3520.get(0);
        mod_5635.put(47, t);
    endrule
    rule rule_126;
        ChannelMessage t;
        t <- mod_5634.get(1);
        mod_44.put(0, t);
    endrule
    rule rule_127;
        ChannelMessage t;
        t <- mod_5634.get(67);
        mod_2948.put(0, t);
    endrule
    rule rule_128;
        ChannelMessage t;
        t <- mod_2068.get(0);
        mod_5635.put(80, t);
    endrule
    rule rule_129;
        ChannelMessage t;
        t <- mod_5633.get(18);
        mod_792.put(1, t);
    endrule
    rule rule_130;
        ChannelMessage t;
        t <- mod_5633.get(84);
        mod_3696.put(1, t);
    endrule
    rule rule_131;
        ChannelMessage t;
        t <- mod_4224.get(0);
        mod_5635.put(31, t);
    endrule
    rule rule_132;
        ChannelMessage t;
        t <- mod_3300.get(0);
        mod_5635.put(52, t);
    endrule
    rule rule_133;
        ChannelMessage t;
        t <- mod_5634.get(82);
        mod_3608.put(0, t);
    endrule
    rule rule_134;
        ChannelMessage t;
        t <- mod_5634.get(95);
        mod_4180.put(0, t);
    endrule
    rule rule_135;
        ChannelMessage t;
        t <- mod_2860.get(0);
        mod_5635.put(62, t);
    endrule
    rule rule_136;
        ChannelMessage t;
        t <- mod_4488.get(0);
        mod_5635.put(25, t);
    endrule
    rule rule_137;
        ChannelMessage t;
        t <- mod_1100.get(0);
        mod_5635.put(102, t);
    endrule
    rule rule_138;
        ChannelMessage t;
        t <- mod_5633.get(5);
        mod_220.put(1, t);
    endrule
    rule rule_139;
        ChannelMessage t;
        t <- mod_5280.get(0);
        mod_5635.put(7, t);
    endrule
    rule rule_140;
        ChannelMessage t;
        t <- mod_4708.get(0);
        mod_5635.put(20, t);
    endrule
    rule rule_141;
        ChannelMessage t;
        t <- mod_4004.get(0);
        mod_5635.put(36, t);
    endrule
    rule rule_142;
        ChannelMessage t;
        t <- mod_5633.get(89);
        mod_3916.put(1, t);
    endrule
    rule rule_143;
        ChannelMessage t;
        t <- mod_5634.get(92);
        mod_4048.put(0, t);
    endrule
    rule rule_144;
        ChannelMessage t;
        t <- mod_792.get(0);
        mod_5635.put(109, t);
    endrule
    rule rule_145;
        ChannelMessage t;
        t <- mod_5634.get(99);
        mod_4356.put(0, t);
    endrule
    rule rule_146;
        ChannelMessage t;
        t <- mod_88.get(0);
        mod_5635.put(125, t);
    endrule
    rule rule_147;
        ChannelMessage t;
        t <- mod_5588.get(0);
        mod_5635.put(0, t);
    endrule
    rule rule_148;
        ChannelMessage t;
        t <- mod_5633.get(57);
        mod_2508.put(1, t);
    endrule
    rule rule_149;
        ChannelMessage t;
        t <- mod_5060.get(0);
        mod_5635.put(12, t);
    endrule
    rule rule_150;
        ChannelMessage t;
        t <- mod_5633.get(121);
        mod_5324.put(1, t);
    endrule
    rule rule_151;
        ChannelMessage t;
        t <- mod_5634.get(59);
        mod_2596.put(0, t);
    endrule
    rule rule_152;
        ChannelMessage t;
        t <- mod_5634.get(98);
        mod_4312.put(0, t);
    endrule
    rule rule_153;
        ChannelMessage t;
        t <- mod_5633.get(47);
        mod_2068.put(1, t);
    endrule
    rule rule_154;
        ChannelMessage t;
        t <- mod_5634.get(14);
        mod_616.put(0, t);
    endrule
    rule rule_155;
        ChannelMessage t;
        t <- mod_5633.get(106);
        mod_4664.put(1, t);
    endrule
    rule rule_156;
        ChannelMessage t;
        t <- mod_3476.get(0);
        mod_5635.put(48, t);
    endrule
    rule rule_157;
        ChannelMessage t;
        t <- mod_4136.get(0);
        mod_5635.put(33, t);
    endrule
    rule rule_158;
        ChannelMessage t;
        t <- mod_5634.get(44);
        mod_1936.put(0, t);
    endrule
    rule rule_159;
        ChannelMessage t;
        t <- mod_5633.get(88);
        mod_3872.put(1, t);
    endrule
    rule rule_160;
        ChannelMessage t;
        t <- mod_4620.get(0);
        mod_5635.put(22, t);
    endrule
    rule rule_161;
        ChannelMessage t;
        t <- mod_5633.get(6);
        mod_264.put(1, t);
    endrule
    rule rule_162;
        ChannelMessage t;
        t <- mod_5633.get(24);
        mod_1056.put(1, t);
    endrule
    rule rule_163;
        ChannelMessage t;
        t <- mod_5633.get(23);
        mod_1012.put(1, t);
    endrule
    rule rule_164;
        ChannelMessage t;
        t <- mod_5633.get(32);
        mod_1408.put(1, t);
    endrule
    rule rule_165;
        ChannelMessage t;
        t <- mod_5633.get(40);
        mod_1760.put(1, t);
    endrule
    rule rule_166;
        ChannelMessage t;
        t <- mod_5633.get(114);
        mod_5016.put(1, t);
    endrule
    rule rule_167;
        ChannelMessage t;
        t <- mod_2508.get(0);
        mod_5635.put(70, t);
    endrule
    rule rule_168;
        ChannelMessage t;
        t <- mod_5633.get(42);
        mod_1848.put(1, t);
    endrule
    rule rule_169;
        ChannelMessage t;
        t <- mod_5634.get(19);
        mod_836.put(0, t);
    endrule
    rule rule_170;
        ChannelMessage t;
        t <- mod_5634.get(20);
        mod_880.put(0, t);
    endrule
    rule rule_171;
        ChannelMessage t;
        t <- mod_5634.get(35);
        mod_1540.put(0, t);
    endrule
    rule rule_172;
        ChannelMessage t;
        t <- mod_5633.get(99);
        mod_4356.put(1, t);
    endrule
    rule rule_173;
        ChannelMessage t;
        t <- mod_5633.get(16);
        mod_704.put(1, t);
    endrule
    rule rule_174;
        ChannelMessage t;
        t <- mod_5634.get(53);
        mod_2332.put(0, t);
    endrule
    rule rule_175;
        ChannelMessage t;
        t <- mod_5634.get(56);
        mod_2464.put(0, t);
    endrule
    rule rule_176;
        ChannelMessage t;
        t <- mod_616.get(0);
        mod_5635.put(113, t);
    endrule
    rule rule_177;
        ChannelMessage t;
        t <- mod_1848.get(0);
        mod_5635.put(85, t);
    endrule
    rule rule_178;
        ChannelMessage t;
        t <- mod_5633.get(60);
        mod_2640.put(1, t);
    endrule
    rule rule_179;
        ChannelMessage t;
        t <- mod_5634.get(3);
        mod_132.put(0, t);
    endrule
    rule rule_180;
        ChannelMessage t;
        t <- mod_5634.get(5);
        mod_220.put(0, t);
    endrule
    rule rule_181;
        ChannelMessage t;
        t <- mod_5634.get(52);
        mod_2288.put(0, t);
    endrule
    rule rule_182;
        ChannelMessage t;
        t <- mod_5634.get(57);
        mod_2508.put(0, t);
    endrule
    rule rule_183;
        ChannelMessage t;
        t <- mod_2728.get(0);
        mod_5635.put(65, t);
    endrule
    rule rule_184;
        ChannelMessage t;
        t <- mod_5634.get(65);
        mod_2860.put(0, t);
    endrule
    rule rule_185;
        ChannelMessage t;
        t <- mod_5633.get(90);
        mod_3960.put(1, t);
    endrule
    rule rule_186;
        ChannelMessage t;
        t <- mod_1408.get(0);
        mod_5635.put(95, t);
    endrule
    rule rule_187;
        ChannelMessage t;
        t <- mod_5633.get(91);
        mod_4004.put(1, t);
    endrule
    rule rule_188;
        ChannelMessage t;
        t <- mod_5634.get(36);
        mod_1584.put(0, t);
    endrule
    rule rule_189;
        ChannelMessage t;
        t <- mod_5192.get(0);
        mod_5635.put(9, t);
    endrule
    rule rule_190;
        ChannelMessage t;
        t <- mod_5633.get(124);
        mod_5456.put(1, t);
    endrule
    rule rule_191;
        ChannelMessage t;
        t <- mod_1584.get(0);
        mod_5635.put(91, t);
    endrule
    rule rule_192;
        ChannelMessage t;
        t <- mod_5634.get(69);
        mod_3036.put(0, t);
    endrule
    rule rule_193;
        ChannelMessage t;
        t <- mod_5634.get(2);
        mod_88.put(0, t);
    endrule
    rule rule_194;
        ChannelMessage t;
        t <- mod_5634.get(91);
        mod_4004.put(0, t);
    endrule
    rule rule_195;
        ChannelMessage t;
        t <- mod_5634.get(51);
        mod_2244.put(0, t);
    endrule
    rule rule_196;
        ChannelMessage t;
        t <- mod_4180.get(0);
        mod_5635.put(32, t);
    endrule
    rule rule_197;
        ChannelMessage t;
        t <- mod_5636.get(0);
        mod_5634.put(0, t);
    endrule
    rule rule_198;
        ChannelMessage t;
        t <- mod_5634.get(27);
        mod_1188.put(0, t);
    endrule
    rule rule_199;
        ChannelMessage t;
        t <- mod_5634.get(70);
        mod_3080.put(0, t);
    endrule
    rule rule_200;
        ChannelMessage t;
        t <- mod_5643.get(0);
        mod_5634.put(1, t);
    endrule
    rule rule_201;
        ChannelMessage t;
        t <- mod_5634.get(41);
        mod_1804.put(0, t);
    endrule
    rule rule_202;
        ChannelMessage t;
        t <- mod_5633.get(35);
        mod_1540.put(1, t);
    endrule
    rule rule_203;
        ChannelMessage t;
        t <- mod_5634.get(58);
        mod_2552.put(0, t);
    endrule
    rule rule_204;
        ChannelMessage t;
        t <- mod_5634.get(111);
        mod_4884.put(0, t);
    endrule
    rule rule_205;
        ChannelMessage t;
        t <- mod_5633.get(22);
        mod_968.put(1, t);
    endrule
    rule rule_206;
        ChannelMessage t;
        t <- mod_5634.get(4);
        mod_176.put(0, t);
    endrule
    rule rule_207;
        ChannelMessage t;
        t <- mod_5634.get(97);
        mod_4268.put(0, t);
    endrule
    rule rule_208;
        ChannelMessage t;
        t <- mod_5633.get(17);
        mod_748.put(1, t);
    endrule
    rule rule_209;
        ChannelMessage t;
        t <- mod_5633.get(34);
        mod_1496.put(1, t);
    endrule
    rule rule_210;
        ChannelMessage t;
        t <- mod_5633.get(14);
        mod_616.put(1, t);
    endrule
    rule rule_211;
        ChannelMessage t;
        t <- mod_5633.get(43);
        mod_1892.put(1, t);
    endrule
    rule rule_212;
        ChannelMessage t;
        t <- mod_5633.get(126);
        mod_5544.put(1, t);
    endrule
    rule rule_213;
        ChannelMessage t;
        t <- mod_5634.get(21);
        mod_924.put(0, t);
    endrule
    rule rule_214;
        ChannelMessage t;
        t <- mod_5634.get(33);
        mod_1452.put(0, t);
    endrule
    rule rule_215;
        ChannelMessage t;
        t <- mod_3344.get(0);
        mod_5635.put(51, t);
    endrule
    rule rule_216;
        ChannelMessage t;
        t <- mod_5633.get(74);
        mod_3256.put(1, t);
    endrule
    rule rule_217;
        ChannelMessage t;
        t <- mod_5633.get(120);
        mod_5280.put(1, t);
    endrule
    rule rule_218;
        ChannelMessage t;
        t <- mod_5633.get(33);
        mod_1452.put(1, t);
    endrule
    rule rule_219;
        ChannelMessage t;
        t <- mod_5634.get(96);
        mod_4224.put(0, t);
    endrule
    rule rule_220;
        ChannelMessage t;
        t <- mod_5633.get(66);
        mod_2904.put(1, t);
    endrule
    rule rule_221;
        ChannelMessage t;
        t <- mod_5634.get(102);
        mod_4488.put(0, t);
    endrule
    rule rule_222;
        ChannelMessage t;
        t <- mod_5634.get(108);
        mod_4752.put(0, t);
    endrule
    rule rule_223;
        ChannelMessage t;
        t <- mod_5639.get(0);
        mod_5633.put(1, t);
    endrule
    rule rule_224;
        ChannelMessage t;
        t <- mod_5633.get(10);
        mod_440.put(1, t);
    endrule
    rule rule_225;
        ChannelMessage t;
        t <- mod_5647.get(0);
        mod_5643.put(0, t);
    endrule
    rule rule_226;
        ChannelMessage t;
        t <- mod_1496.get(0);
        mod_5635.put(93, t);
    endrule
    rule rule_227;
        ChannelMessage t;
        t <- mod_5633.get(79);
        mod_3476.put(1, t);
    endrule
    rule rule_228;
        ChannelMessage t;
        t <- mod_5633.get(94);
        mod_4136.put(1, t);
    endrule
    rule rule_229;
        ChannelMessage t;
        t <- mod_3168.get(0);
        mod_5635.put(55, t);
    endrule
    rule rule_230;
        ChannelMessage t;
        t <- mod_5645.get(0);
        mod_5638.put(0, t);
    endrule
    rule rule_231;
        ChannelMessage t;
        t <- mod_572.get(0);
        mod_5635.put(114, t);
    endrule
    rule rule_232;
        ChannelMessage t;
        t <- mod_5634.get(84);
        mod_3696.put(0, t);
    endrule
    rule rule_233;
        ChannelMessage t;
        t <- mod_3212.get(0);
        mod_5635.put(54, t);
    endrule
    rule rule_234;
        ChannelMessage t;
        t <- mod_5633.get(69);
        mod_3036.put(1, t);
    endrule
    rule rule_235;
        ChannelMessage t;
        t <- mod_5634.get(80);
        mod_3520.put(0, t);
    endrule
    rule rule_236;
        ChannelMessage t;
        t <- mod_0.get(0);
        mod_5635.put(127, t);
    endrule
    rule rule_237;
        ChannelMessage t;
        t <- mod_5633.get(100);
        mod_4400.put(1, t);
    endrule
    rule rule_238;
        ChannelMessage t;
        t <- mod_5634.get(17);
        mod_748.put(0, t);
    endrule
    rule rule_239;
        ChannelMessage t;
        t <- mod_3124.get(0);
        mod_5635.put(56, t);
    endrule
    rule rule_240;
        ChannelMessage t;
        t <- mod_5634.get(42);
        mod_1848.put(0, t);
    endrule
    rule rule_241;
        ChannelMessage t;
        t <- mod_5634.get(79);
        mod_3476.put(0, t);
    endrule
    rule rule_242;
        ChannelMessage t;
        t <- mod_1716.get(0);
        mod_5635.put(88, t);
    endrule
    rule rule_243;
        ChannelMessage t;
        t <- mod_5633.get(1);
        mod_44.put(1, t);
    endrule
    rule rule_244;
        ChannelMessage t;
        t <- mod_5634.get(12);
        mod_528.put(0, t);
    endrule
    rule rule_245;
        ChannelMessage t;
        t <- mod_5633.get(8);
        mod_352.put(1, t);
    endrule
    rule rule_246;
        ChannelMessage t;
        t <- mod_924.get(0);
        mod_5635.put(106, t);
    endrule
    rule rule_247;
        ChannelMessage t;
        t <- mod_5633.get(104);
        mod_4576.put(1, t);
    endrule
    rule rule_248;
        ChannelMessage t;
        t <- mod_5634.get(119);
        mod_5236.put(0, t);
    endrule
    rule rule_249;
        ChannelMessage t;
        t <- mod_5634.get(120);
        mod_5280.put(0, t);
    endrule
    rule rule_250;
        ChannelMessage t;
        t <- mod_5633.get(98);
        mod_4312.put(1, t);
    endrule
    rule rule_251;
        ChannelMessage t;
        t <- mod_4664.get(0);
        mod_5635.put(21, t);
    endrule
    rule rule_252;
        ChannelMessage t;
        t <- mod_5634.get(24);
        mod_1056.put(0, t);
    endrule
    rule rule_253;
        ChannelMessage t;
        t <- mod_5634.get(40);
        mod_1760.put(0, t);
    endrule
    rule rule_254;
        ChannelMessage t;
        t <- mod_5634.get(63);
        mod_2772.put(0, t);
    endrule
    rule rule_255;
        ChannelMessage t;
        t <- mod_5633.get(76);
        mod_3344.put(1, t);
    endrule
    rule rule_256;
        ChannelMessage t;
        t <- mod_5634.get(86);
        mod_3784.put(0, t);
    endrule
    rule rule_257;
        ChannelMessage t;
        t <- mod_5634.get(37);
        mod_1628.put(0, t);
    endrule
    rule rule_258;
        ChannelMessage t;
        t <- mod_5634.get(48);
        mod_2112.put(0, t);
    endrule
    rule rule_259;
        ChannelMessage t;
        t <- mod_5634.get(78);
        mod_3432.put(0, t);
    endrule
    rule rule_260;
        ChannelMessage t;
        t <- mod_5646.get(0);
        mod_5635.put(128, t);
    endrule
    rule rule_261;
        ChannelMessage t;
        t <- mod_5638.get(0);
        mod_5638.put(1, t);
    endrule
    rule rule_262;
        ChannelMessage t;
        t <- mod_5633.get(109);
        mod_4796.put(1, t);
    endrule
    rule rule_263;
        ChannelMessage t;
        t <- mod_132.get(0);
        mod_5635.put(124, t);
    endrule
    rule rule_264;
        ChannelMessage t;
        t <- mod_5635.get(0);
        mod_5645.put(0, t);
    endrule
    rule rule_265;
        ChannelMessage t;
        t <- mod_5634.get(46);
        mod_2024.put(0, t);
    endrule
    rule rule_266;
        ChannelMessage t;
        t <- mod_5633.get(85);
        mod_3740.put(1, t);
    endrule
    rule rule_267;
        ChannelMessage t;
        t <- mod_5634.get(50);
        mod_2200.put(0, t);
    endrule
    rule rule_268;
        ChannelMessage t;
        t <- mod_1452.get(0);
        mod_5635.put(94, t);
    endrule
    rule rule_269;
        ChannelMessage t;
        t <- mod_5633.get(27);
        mod_1188.put(1, t);
    endrule
    rule rule_270;
        ChannelMessage t;
        t <- mod_5634.get(105);
        mod_4620.put(0, t);
    endrule
    rule rule_271;
        ChannelMessage t;
        t <- mod_5634.get(23);
        mod_1012.put(0, t);
    endrule
    rule rule_272;
        ChannelMessage t;
        t <- mod_5634.get(55);
        mod_2420.put(0, t);
    endrule
    rule rule_273;
        ChannelMessage t;
        t <- mod_3784.get(0);
        mod_5635.put(41, t);
    endrule
    rule rule_274;
        ChannelMessage t;
        t <- mod_3960.get(0);
        mod_5635.put(37, t);
    endrule
    rule rule_275;
        ChannelMessage t;
        t <- mod_2244.get(0);
        mod_5635.put(76, t);
    endrule
    rule rule_276;
        ChannelMessage t;
        t <- mod_5633.get(116);
        mod_5104.put(1, t);
    endrule
    rule rule_277;
        ChannelMessage t;
        t <- mod_5633.get(56);
        mod_2464.put(1, t);
    endrule
    rule rule_278;
        ChannelMessage t;
        t <- mod_5634.get(26);
        mod_1144.put(0, t);
    endrule
    rule rule_279;
        ChannelMessage t;
        t <- mod_5634.get(81);
        mod_3564.put(0, t);
    endrule
    rule rule_280;
        ChannelMessage t;
        t <- mod_5634.get(118);
        mod_5192.put(0, t);
    endrule
    rule rule_281;
        ChannelMessage t;
        t <- mod_5633.get(39);
        mod_1716.put(1, t);
    endrule
    rule rule_282;
        ChannelMessage t;
        t <- mod_5634.get(45);
        mod_1980.put(0, t);
    endrule
    rule rule_283;
        ChannelMessage t;
        t <- mod_220.get(0);
        mod_5635.put(122, t);
    endrule
    rule rule_284;
        ChannelMessage t;
        t <- mod_1672.get(0);
        mod_5635.put(89, t);
    endrule
    rule rule_285;
        ChannelMessage t;
        t <- mod_2464.get(0);
        mod_5635.put(71, t);
    endrule
    rule rule_286;
        ChannelMessage t;
        t <- mod_5368.get(0);
        mod_5635.put(5, t);
    endrule
    rule rule_287;
        ChannelMessage t;
        t <- mod_5634.get(34);
        mod_1496.put(0, t);
    endrule
    rule rule_288;
        ChannelMessage t;
        t <- mod_5633.get(45);
        mod_1980.put(1, t);
    endrule
    rule rule_289;
        ChannelMessage t;
        t <- mod_5633.get(77);
        mod_3388.put(1, t);
    endrule
    rule rule_290;
        ChannelMessage t;
        t <- mod_3652.get(0);
        mod_5635.put(44, t);
    endrule
    rule rule_291;
        ChannelMessage t;
        t <- mod_5633.get(2);
        mod_88.put(1, t);
    endrule
    rule rule_292;
        ChannelMessage t;
        t <- mod_5633.get(4);
        mod_176.put(1, t);
    endrule
    rule rule_293;
        ChannelMessage t;
        t <- mod_704.get(0);
        mod_5635.put(111, t);
    endrule
    rule rule_294;
        ChannelMessage t;
        t <- mod_2552.get(0);
        mod_5635.put(69, t);
    endrule
    rule rule_295;
        ChannelMessage t;
        t <- mod_5633.get(52);
        mod_2288.put(1, t);
    endrule
    rule rule_296;
        ChannelMessage t;
        t <- mod_5633.get(107);
        mod_4708.put(1, t);
    endrule
    rule rule_297;
        ChannelMessage t;
        t <- mod_5633.get(123);
        mod_5412.put(1, t);
    endrule
    rule rule_298;
        ChannelMessage t;
        t <- mod_5633.get(9);
        mod_396.put(1, t);
    endrule
    rule rule_299;
        ChannelMessage t;
        t <- mod_1012.get(0);
        mod_5635.put(104, t);
    endrule
    rule rule_300;
        ChannelMessage t;
        t <- mod_5148.get(0);
        mod_5635.put(10, t);
    endrule
    rule rule_301;
        ChannelMessage t;
        t <- mod_5634.get(11);
        mod_484.put(0, t);
    endrule
    rule rule_302;
        ChannelMessage t;
        t <- mod_5633.get(119);
        mod_5236.put(1, t);
    endrule
    rule rule_303;
        ChannelMessage t;
        t <- mod_5634.get(87);
        mod_3828.put(0, t);
    endrule
    rule rule_304;
        ChannelMessage t;
        t <- mod_5633.get(26);
        mod_1144.put(1, t);
    endrule
    rule rule_305;
        ChannelMessage t;
        t <- mod_5634.get(112);
        mod_4928.put(0, t);
    endrule
    rule rule_306;
        ChannelMessage t;
        t <- mod_5634.get(113);
        mod_4972.put(0, t);
    endrule
    rule rule_307;
        ChannelMessage t;
        t <- mod_4576.get(0);
        mod_5635.put(23, t);
    endrule
    rule rule_308;
        ChannelMessage t;
        t <- mod_5633.get(54);
        mod_2376.put(1, t);
    endrule
    rule rule_309;
        ChannelMessage t;
        t <- mod_4884.get(0);
        mod_5635.put(16, t);
    endrule
    rule rule_310;
        ChannelMessage t;
        t <- mod_5634.get(116);
        mod_5104.put(0, t);
    endrule
    rule rule_311;
        ChannelMessage t;
        t <- mod_5456.get(0);
        mod_5635.put(3, t);
    endrule
    rule rule_312;
        ChannelMessage t;
        t <- mod_5648.get(0);
        mod_5639.put(0, t);
    endrule
    rule rule_313;
        ChannelMessage t;
        t <- mod_1276.get(0);
        mod_5635.put(98, t);
    endrule
    rule rule_314;
        ChannelMessage t;
        t <- mod_5633.get(97);
        mod_4268.put(1, t);
    endrule
    rule rule_315;
        ChannelMessage t;
        t <- mod_5634.get(61);
        mod_2684.put(0, t);
    endrule
    rule rule_316;
        ChannelMessage t;
        t <- mod_748.get(0);
        mod_5635.put(110, t);
    endrule
    rule rule_317;
        ChannelMessage t;
        t <- mod_3872.get(0);
        mod_5635.put(39, t);
    endrule
    rule rule_318;
        ChannelMessage t;
        t <- mod_5634.get(13);
        mod_572.put(0, t);
    endrule
    rule rule_319;
        ChannelMessage t;
        t <- mod_2816.get(0);
        mod_5635.put(63, t);
    endrule
    rule rule_320;
        ChannelMessage t;
        t <- mod_5634.get(73);
        mod_3212.put(0, t);
    endrule
    rule rule_321;
        ChannelMessage t;
        t <- mod_1980.get(0);
        mod_5635.put(82, t);
    endrule
    rule rule_322;
        ChannelMessage t;
        t <- mod_5634.get(125);
        mod_5500.put(0, t);
    endrule
    rule rule_323;
        ChannelMessage t;
        t <- mod_5633.get(108);
        mod_4752.put(1, t);
    endrule
    rule rule_324;
        ChannelMessage t;
        t <- mod_5634.get(43);
        mod_1892.put(0, t);
    endrule
    rule rule_325;
        ChannelMessage t;
        t <- mod_5324.get(0);
        mod_5635.put(6, t);
    endrule
    rule rule_326;
        ChannelMessage t;
        t <- mod_2684.get(0);
        mod_5635.put(66, t);
    endrule
    rule rule_327;
        ChannelMessage t;
        t <- mod_5104.get(0);
        mod_5635.put(11, t);
    endrule
    rule rule_328;
        ChannelMessage t;
        t <- mod_5634.get(15);
        mod_660.put(0, t);
    endrule
    rule rule_329;
        ChannelMessage t;
        t <- mod_4972.get(0);
        mod_5635.put(14, t);
    endrule
    rule rule_330;
        ChannelMessage t;
        t <- mod_1892.get(0);
        mod_5635.put(84, t);
    endrule
    rule rule_331;
        ChannelMessage t;
        t <- mod_1144.get(0);
        mod_5635.put(101, t);
    endrule
    rule rule_332;
        ChannelMessage t;
        t <- mod_5634.get(123);
        mod_5412.put(0, t);
    endrule
    rule rule_333;
        ChannelMessage t;
        t <- mod_5633.get(65);
        mod_2860.put(1, t);
    endrule
    rule rule_334;
        ChannelMessage t;
        t <- mod_5633.get(30);
        mod_1320.put(1, t);
    endrule
    rule rule_335;
        ChannelMessage t;
        t <- mod_396.get(0);
        mod_5635.put(118, t);
    endrule
    rule rule_336;
        ChannelMessage t;
        t <- mod_5634.get(8);
        mod_352.put(0, t);
    endrule
    rule rule_337;
        ChannelMessage t;
        t <- mod_5633.get(59);
        mod_2596.put(1, t);
    endrule
    rule rule_338;
        ChannelMessage t;
        t <- mod_5634.get(75);
        mod_3300.put(0, t);
    endrule
    rule rule_339;
        ChannelMessage t;
        t <- mod_5633.get(83);
        mod_3652.put(1, t);
    endrule
    rule rule_340;
        ChannelMessage t;
        t <- mod_5634.get(77);
        mod_3388.put(0, t);
    endrule
    rule rule_341;
        ChannelMessage t;
        t <- mod_5016.get(0);
        mod_5635.put(13, t);
    endrule
    rule rule_342;
        ChannelMessage t;
        t <- mod_5633.get(67);
        mod_2948.put(1, t);
    endrule
    rule rule_343;
        ChannelMessage t;
        t <- mod_5634.get(100);
        mod_4400.put(0, t);
    endrule
    rule rule_344;
        ChannelMessage t;
        t <- mod_44.get(0);
        mod_5635.put(126, t);
    endrule
    rule rule_345;
        ChannelMessage t;
        t <- mod_5634.get(124);
        mod_5456.put(0, t);
    endrule
    rule rule_346;
        ChannelMessage t;
        t <- mod_1232.get(0);
        mod_5635.put(99, t);
    endrule
    rule rule_347;
        ChannelMessage t;
        t <- mod_5633.get(93);
        mod_4092.put(1, t);
    endrule
    rule rule_348;
        ChannelMessage t;
        t <- mod_5640.get(0);
        mod_5646.put(0, t);
    endrule
    rule rule_349;
        ChannelMessage t;
        t <- mod_440.get(0);
        mod_5635.put(117, t);
    endrule
    rule rule_350;
        ChannelMessage t;
        t <- mod_5634.get(76);
        mod_3344.put(0, t);
    endrule
    rule rule_351;
        ChannelMessage t;
        t <- mod_5633.get(38);
        mod_1672.put(1, t);
    endrule
    rule rule_352;
        ChannelMessage t;
        t <- mod_5634.get(83);
        mod_3652.put(0, t);
    endrule
    rule rule_353;
        ChannelMessage t;
        t <- mod_4928.get(0);
        mod_5635.put(15, t);
    endrule
    rule rule_354;
        ChannelMessage t;
        t <- mod_5634.get(71);
        mod_3124.put(0, t);
    endrule
    rule rule_355;
        ChannelMessage t;
        t <- mod_5634.get(101);
        mod_4444.put(0, t);
    endrule
    rule rule_356;
        ChannelMessage t;
        t <- mod_352.get(0);
        mod_5635.put(119, t);
    endrule
    rule rule_357;
        ChannelMessage t;
        t <- mod_5634.get(104);
        mod_4576.put(0, t);
    endrule
    rule rule_358;
        ChannelMessage t;
        t <- mod_5633.get(125);
        mod_5500.put(1, t);
    endrule
    rule rule_359;
        ChannelMessage t;
        t <- mod_5634.get(122);
        mod_5368.put(0, t);
    endrule
    rule rule_360;
        ChannelMessage t;
        t <- mod_5634.get(126);
        mod_5544.put(0, t);
    endrule
    rule rule_361;
        ChannelMessage t;
        t <- mod_5644.get(0);
        mod_5633.put(0, t);
    endrule
    rule rule_362;
        ChannelMessage t;
        t <- mod_3080.get(0);
        mod_5635.put(57, t);
    endrule
    rule rule_363;
        ChannelMessage t;
        t <- mod_5633.get(3);
        mod_132.put(1, t);
    endrule
    rule rule_364;
        ChannelMessage t;
        t <- mod_5634.get(9);
        mod_396.put(0, t);
    endrule
    rule rule_365;
        ChannelMessage t;
        t <- mod_5634.get(38);
        mod_1672.put(0, t);
    endrule
    rule rule_366;
        ChannelMessage t;
        t <- mod_2948.get(0);
        mod_5635.put(60, t);
    endrule
    rule rule_367;
        ChannelMessage t;
        t <- mod_5633.get(46);
        mod_2024.put(1, t);
    endrule
    rule rule_368;
        ChannelMessage t;
        t <- mod_5500.get(0);
        mod_5635.put(2, t);
    endrule
    rule rule_369;
        ChannelMessage t;
        t <- mod_4840.get(0);
        mod_5635.put(17, t);
    endrule
    rule rule_370;
        ChannelMessage t;
        t <- mod_5634.get(39);
        mod_1716.put(0, t);
    endrule
    rule rule_371;
        ChannelMessage t;
        t <- mod_5634.get(88);
        mod_3872.put(0, t);
    endrule
    rule rule_372;
        ChannelMessage t;
        t <- mod_5634.get(110);
        mod_4840.put(0, t);
    endrule
    rule rule_373;
        ChannelMessage t;
        t <- mod_5634.get(90);
        mod_3960.put(0, t);
    endrule
    rule rule_374;
        ChannelMessage t;
        t <- mod_5633.get(29);
        mod_1276.put(1, t);
    endrule
    rule rule_375;
        ChannelMessage t;
        t <- mod_5633.get(87);
        mod_3828.put(1, t);
    endrule
    rule rule_376;
        ChannelMessage t;
        t <- mod_660.get(0);
        mod_5635.put(112, t);
    endrule
    rule rule_377;
        ChannelMessage t;
        t <- mod_3388.get(0);
        mod_5635.put(50, t);
    endrule
    rule rule_378;
        ChannelMessage t;
        t <- mod_5412.get(0);
        mod_5635.put(4, t);
    endrule
    rule rule_379;
        ChannelMessage t;
        t <- mod_2772.get(0);
        mod_5635.put(64, t);
    endrule
    rule rule_380;
        ChannelMessage t;
        t <- mod_4444.get(0);
        mod_5635.put(26, t);
    endrule
    rule rule_381;
        ChannelMessage t;
        t <- mod_5633.get(61);
        mod_2684.put(1, t);
    endrule
    rule rule_382;
        ChannelMessage t;
        t <- mod_5633.get(11);
        mod_484.put(1, t);
    endrule
    rule rule_383;
        ChannelMessage t;
        t <- mod_4752.get(0);
        mod_5635.put(19, t);
    endrule
    rule rule_384;
        ChannelMessage t;
        t <- mod_1760.get(0);
        mod_5635.put(87, t);
    endrule
    rule rule_385;
        ChannelMessage t;
        t <- mod_5633.get(101);
        mod_4444.put(1, t);
    endrule
    rule rule_386;
        ChannelMessage t;
        t <- mod_880.get(0);
        mod_5635.put(107, t);
    endrule
    rule rule_387;
        ChannelMessage t;
        t <- mod_1936.get(0);
        mod_5635.put(83, t);
    endrule
    rule rule_388;
        ChannelMessage t;
        t <- mod_5634.get(6);
        mod_264.put(0, t);
    endrule
    rule rule_389;
        ChannelMessage t;
        t <- mod_4092.get(0);
        mod_5635.put(34, t);
    endrule
    rule rule_390;
        ChannelMessage t;
        t <- mod_5633.get(41);
        mod_1804.put(1, t);
    endrule
    rule rule_391;
        ChannelMessage t;
        t <- mod_5634.get(32);
        mod_1408.put(0, t);
    endrule
    rule rule_392;
        ChannelMessage t;
        t <- mod_5634.get(121);
        mod_5324.put(0, t);
    endrule
    rule rule_393;
        ChannelMessage t;
        t <- mod_1364.get(0);
        mod_5635.put(96, t);
    endrule
    rule rule_394;
        ChannelMessage t;
        t <- mod_5633.get(81);
        mod_3564.put(1, t);
    endrule
    rule rule_395;
        ChannelMessage t;
        t <- mod_5634.get(29);
        mod_1276.put(0, t);
    endrule
    rule rule_396;
        ChannelMessage t;
        t <- mod_1540.get(0);
        mod_5635.put(92, t);
    endrule
    rule rule_397;
        ChannelMessage t;
        t <- mod_5633.get(44);
        mod_1936.put(1, t);
    endrule
    rule rule_398;
        ChannelMessage t;
        t <- mod_5634.get(89);
        mod_3916.put(0, t);
    endrule
    rule rule_399;
        ChannelMessage t;
        t <- mod_5633.get(117);
        mod_5148.put(1, t);
    endrule
    rule rule_400;
        ChannelMessage t;
        t <- mod_4268.get(0);
        mod_5635.put(30, t);
    endrule

endmodule
endpackage
